--2020-02-25 22:13:57--  http://libroslibres.uls.edu.sv/politica/militares_junto_al_pueblo.pdf%0D
Resolving libroslibres.uls.edu.sv (libroslibres.uls.edu.sv)... 72.249.68.209
Connecting to libroslibres.uls.edu.sv (libroslibres.uls.edu.sv)|72.249.68.209|:80... failed: Connection timed out.
Giving up.

--2020-02-25 22:14:23--  http://libroslibres.uls.edu.sv/politica/militares_junto_al_pueblo.pdf%0D
Resolving libroslibres.uls.edu.sv (libroslibres.uls.edu.sv)... 72.249.68.209
Connecting to libroslibres.uls.edu.sv (libroslibres.uls.edu.sv)|72.249.68.209|:80... failed: Connection timed out.
Giving up.

