--2020-03-02 03:24:18--  http://www.jurisprudencia.gob.sv/publicados/Juris_Publicados_Junio2019v3.pdf
Resolving www.jurisprudencia.gob.sv (www.jurisprudencia.gob.sv)... 200.31.169.67
Connecting to www.jurisprudencia.gob.sv (www.jurisprudencia.gob.sv)|200.31.169.67|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 1504544 (1.4M) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  3%  766K 15s
    50K .......... .......... .......... .......... ..........  6% 3.01M 9s
   100K .......... .......... .......... .......... .......... 10%  125M 6s
   150K .......... .......... .......... .......... .......... 13% 3.16M 5s
   200K .......... .......... .......... .......... .......... 17% 54.4M 4s
   250K .......... .......... .......... .......... .......... 20%  275M 3s
   300K .......... .......... .......... .......... .......... 23% 3.26M 3s
   350K .......... .......... .......... .......... .......... 27% 74.4M 3s
   400K .......... .......... .......... .......... .......... 30%  105M 2s
   450K .......... .......... .......... .......... .......... 34% 3.38M 2s
   500K .......... .......... .......... .......... .......... 37% 82.5M 2s
   550K .......... .......... .......... .......... .......... 40%  160M 2s
   600K .......... .......... .......... .......... .......... 44%  124M 1s
   650K .......... .......... .......... .......... .......... 47%  145M 1s
   700K .......... .......... .......... .......... .......... 51% 3.43M 1s
   750K .......... .......... .......... .......... .......... 54%  113M 1s
   800K .......... .......... .......... .......... .......... 57% 94.7M 1s
   850K .......... .......... .......... .......... .......... 61%  238M 1s
   900K .......... .......... .......... .......... .......... 64%  203M 1s
   950K .......... .......... .......... .......... .......... 68%  106M 1s
  1000K .......... .......... .......... .......... .......... 71%  194M 0s
  1050K .......... .......... .......... .......... .......... 74% 3.53M 0s
  1100K .......... .......... .......... .......... .......... 78%  189M 0s
  1150K .......... .......... .......... .......... .......... 81%  102M 0s
  1200K .......... .......... .......... .......... .......... 85%  558M 0s
  1250K .......... .......... .......... .......... .......... 88%  190M 0s
  1300K .......... .......... .......... .......... .......... 91%  136M 0s
  1350K .......... .......... .......... .......... .......... 95%  196M 0s
  1400K .......... .......... .......... .......... .......... 98%  407M 0s
  1450K .......... .........                                  100% 97.1M=1.4s

2020-03-02 03:24:20 (8.90 Mb/s) - ‘/dev/null’ saved [1504544/1504544]

