--2020-03-02 03:26:19--  http://www.promerica.com.sv/media/1229/reglamento.pdf
Resolving www.promerica.com.sv (www.promerica.com.sv)... 45.60.154.167
Connecting to www.promerica.com.sv (www.promerica.com.sv)|45.60.154.167|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: https://www.promerica.com.sv [following]
--2020-03-02 03:26:19--  https://www.promerica.com.sv/
Connecting to www.promerica.com.sv (www.promerica.com.sv)|45.60.154.167|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 1.60M
    50K .......... ....                                        92.9M=0.3s

2020-03-02 03:26:21 (2.06 Mb/s) - ‘/dev/null’ saved [66106]

