--2020-03-02 03:27:11--  http://tienda.movistar.com.sv/tv/Movistar_TvHD_Manual_Uso.pdf
Resolving tienda.movistar.com.sv (tienda.movistar.com.sv)... 72.47.233.224
Connecting to tienda.movistar.com.sv (tienda.movistar.com.sv)|72.47.233.224|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 3520006 (3.4M) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  1% 1.45M 19s
    50K .......... .......... .......... .......... ..........  2% 2.88M 14s
   100K .......... .......... .......... .......... ..........  4% 2.92M 12s
   150K .......... .......... .......... .......... ..........  5% 2.97M 11s
   200K .......... .......... .......... .......... ..........  7%  106M 9s
   250K .......... .......... .......... .......... ..........  8% 2.99M 9s
   300K .......... .......... .......... .......... .......... 10% 96.2M 7s
   350K .......... .......... .......... .......... .......... 11% 86.4M 6s
   400K .......... .......... .......... .......... .......... 13% 3.10M 7s
   450K .......... .......... .......... .......... .......... 14%  220M 6s
   500K .......... .......... .......... .......... .......... 15%  109M 5s
   550K .......... .......... .......... .......... .......... 17% 94.2M 5s
   600K .......... .......... .......... .......... .......... 18% 3.15M 5s
   650K .......... .......... .......... .......... .......... 20% 88.1M 4s
   700K .......... .......... .......... .......... .......... 21%  180M 4s
   750K .......... .......... .......... .......... .......... 23%  445M 4s
   800K .......... .......... .......... .......... .......... 24%  135M 3s
   850K .......... .......... .......... .......... .......... 26% 3.16M 4s
   900K .......... .......... .......... .......... .......... 27%  138M 3s
   950K .......... .......... .......... .......... .......... 29%  126M 3s
  1000K .......... .......... .......... .......... .......... 30%  385M 3s
  1050K .......... .......... .......... .......... .......... 31%  184M 3s
  1100K .......... .......... .......... .......... .......... 33%  102M 3s
  1150K .......... .......... .......... .......... .......... 34%  138M 2s
  1200K .......... .......... .......... .......... .......... 36%  741M 2s
  1250K .......... .......... .......... .......... .......... 37% 3.29M 2s
  1300K .......... .......... .......... .......... .......... 39%  106M 2s
  1350K .......... .......... .......... .......... .......... 40%  123M 2s
  1400K .......... .......... .......... .......... .......... 42%  198M 2s
  1450K .......... .......... .......... .......... .......... 43%  173M 2s
  1500K .......... .......... .......... .......... .......... 45%  126M 2s
  1550K .......... .......... .......... .......... .......... 46%  459M 2s
  1600K .......... .......... .......... .......... .......... 47%  411M 2s
  1650K .......... .......... .......... .......... .......... 49%  208M 1s
  1700K .......... .......... .......... .......... .......... 50%  226M 1s
  1750K .......... .......... .......... .......... .......... 52%  351M 1s
  1800K .......... .......... .......... .......... .......... 53% 3.43M 1s
  1850K .......... .......... .......... .......... .......... 55%  246M 1s
  1900K .......... .......... .......... .......... .......... 56%  161M 1s
  1950K .......... .......... .......... .......... .......... 58%  102M 1s
  2000K .......... .......... .......... .......... .......... 59%  180M 1s
  2050K .......... .......... .......... .......... .......... 61%  215M 1s
  2100K .......... .......... .......... .......... .......... 62%  353M 1s
  2150K .......... .......... .......... .......... .......... 63%  204M 1s
  2200K .......... .......... .......... .......... .......... 65%  160M 1s
  2250K .......... .......... .......... .......... .......... 66% 98.9M 1s
  2300K .......... .......... .......... .......... .......... 68% 1.24G 1s
  2350K .......... .......... .......... .......... .......... 69%  222M 1s
  2400K .......... .......... .......... .......... .......... 71%  196M 1s
  2450K .......... .......... .......... .......... .......... 72%  350M 1s
  2500K .......... .......... .......... .......... .......... 74%  197M 1s
  2550K .......... .......... .......... .......... .......... 75% 3.72M 1s
  2600K .......... .......... .......... .......... .......... 77%  117M 1s
  2650K .......... .......... .......... .......... .......... 78%  181M 0s
  2700K .......... .......... .......... .......... .......... 79%  180M 0s
  2750K .......... .......... .......... .......... .......... 81%  263M 0s
  2800K .......... .......... .......... .......... .......... 82%  315M 0s
  2850K .......... .......... .......... .......... .......... 84%  234M 0s
  2900K .......... .......... .......... .......... .......... 85%  240M 0s
  2950K .......... .......... .......... .......... .......... 87%  180M 0s
  3000K .......... .......... .......... .......... .......... 88%  217M 0s
  3050K .......... .......... .......... .......... .......... 90%  509M 0s
  3100K .......... .......... .......... .......... .......... 91%  194M 0s
  3150K .......... .......... .......... .......... .......... 93%  361M 0s
  3200K .......... .......... .......... .......... .......... 94%  241M 0s
  3250K .......... .......... .......... .......... .......... 95%  212M 0s
  3300K .......... .......... .......... .......... .......... 97%  158M 0s
  3350K .......... .......... .......... .......... .......... 98%  279M 0s
  3400K .......... .......... .......... .......              100%  237M=1.7s

2020-03-02 03:27:13 (16.4 Mb/s) - ‘/dev/null’ saved [3520006/3520006]

