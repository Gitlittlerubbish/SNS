--2020-02-25 22:12:49--  https://www.integral.com.sv/asset/documents/859%0D
Resolving www.integral.com.sv (www.integral.com.sv)... 95.216.241.9
Connecting to www.integral.com.sv (www.integral.com.sv)|95.216.241.9|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 6.06M
    50K .......... .......... .......... ....                  1.16G=0.07s

2020-02-25 22:12:49 (10.2 Mb/s) - ‘/dev/null’ saved [86155]

--2020-02-25 22:12:49--  https://www.integral.com.sv/asset/documents/859%0D
Resolving www.integral.com.sv (www.integral.com.sv)... 95.216.241.9
Connecting to www.integral.com.sv (www.integral.com.sv)|95.216.241.9|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 6.55M
    50K .......... .......... .......... ....                  4.09G=0.06s

2020-02-25 22:12:49 (11.0 Mb/s) - ‘/dev/null’ saved [86155]

--2020-02-25 22:13:26--  https://www.integral.com.sv/asset/documents/859%0D
Resolving www.integral.com.sv (www.integral.com.sv)... 95.216.241.9
Connecting to www.integral.com.sv (www.integral.com.sv)|95.216.241.9|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 13.5M
    50K .......... .......... .......... ....                  2.27G=0.03s

2020-02-25 22:13:26 (22.7 Mb/s) - ‘/dev/null’ saved [86155]

--2020-02-25 22:13:26--  https://www.integral.com.sv/asset/documents/859%0D
Resolving www.integral.com.sv (www.integral.com.sv)... 95.216.241.9
Connecting to www.integral.com.sv (www.integral.com.sv)|95.216.241.9|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 5.95M
    50K .......... .......... .......... ....                  2.66G=0.07s

2020-02-25 22:13:27 (10.0 Mb/s) - ‘/dev/null’ saved [86155]

