--2020-03-02 03:27:16--  http://www.ops.com.sv/pdf/205SESeries-Brochure.pdf
Resolving www.ops.com.sv (www.ops.com.sv)... 192.185.148.211
Connecting to www.ops.com.sv (www.ops.com.sv)|192.185.148.211|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 5766625 (5.5M) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  0% 1.68M 27s
    50K .......... .......... .......... .......... ..........  1% 3.30M 20s
   100K .......... .......... .......... .......... ..........  2%  107M 14s
   150K .......... .......... .......... .......... ..........  3%  176M 10s
   200K .......... .......... .......... .......... ..........  4% 3.40M 11s
   250K .......... .......... .......... .......... ..........  5%  183M 9s
   300K .......... .......... .......... .......... ..........  6% 3.51M 9s
   350K .......... .......... .......... .......... ..........  7%  113M 8s
   400K .......... .......... .......... .......... ..........  7%  527M 7s
   450K .......... .......... .......... .......... ..........  8% 88.2M 6s
   500K .......... .......... .......... .......... ..........  9% 53.0M 6s
   550K .......... .......... .......... .......... .......... 10% 3.78M 6s
   600K .......... .......... .......... .......... .......... 11% 79.2M 6s
   650K .......... .......... .......... .......... .......... 12%  410M 5s
   700K .......... .......... .......... .......... .......... 13%  162M 5s
   750K .......... .......... .......... .......... .......... 14% 37.2M 5s
   800K .......... .......... .......... .......... .......... 15% 4.00M 5s
   850K .......... .......... .......... .......... .......... 15%  171M 5s
   900K .......... .......... .......... .......... .......... 16%  722M 4s
   950K .......... .......... .......... .......... .......... 17%  244M 4s
  1000K .......... .......... .......... .......... .......... 18%  195M 4s
  1050K .......... .......... .......... .......... .......... 19%  200M 4s
  1100K .......... .......... .......... .......... .......... 20% 92.9M 3s
  1150K .......... .......... .......... .......... .......... 21% 59.1M 3s
  1200K .......... .......... .......... .......... .......... 22% 4.02M 3s
  1250K .......... .......... .......... .......... .......... 23%  113M 3s
  1300K .......... .......... .......... .......... .......... 23%  107M 3s
  1350K .......... .......... .......... .......... .......... 24%  432M 3s
  1400K .......... .......... .......... .......... .......... 25%  163M 3s
  1450K .......... .......... .......... .......... .......... 26%  207M 3s
  1500K .......... .......... .......... .......... .......... 27%  332M 3s
  1550K .......... .......... .......... .......... .......... 28% 27.9M 3s
  1600K .......... .......... .......... .......... .......... 29%  171M 2s
  1650K .......... .......... .......... .......... .......... 30%  334M 2s
  1700K .......... .......... .......... .......... .......... 31% 4.53M 2s
  1750K .......... .......... .......... .......... .......... 31%  139M 2s
  1800K .......... .......... .......... .......... .......... 32%  291M 2s
  1850K .......... .......... .......... .......... .......... 33%  508M 2s
  1900K .......... .......... .......... .......... .......... 34%  223M 2s
  1950K .......... .......... .......... .......... .......... 35%  395M 2s
  2000K .......... .......... .......... .......... .......... 36%  232M 2s
  2050K .......... .......... .......... .......... .......... 37%  291M 2s
  2100K .......... .......... .......... .......... .......... 38%  563M 2s
  2150K .......... .......... .......... .......... .......... 39%  178M 2s
  2200K .......... .......... .......... .......... .......... 39%  400M 2s
  2250K .......... .......... .......... .......... .......... 40%  207M 2s
  2300K .......... .......... .......... .......... .......... 41%  389M 2s
  2350K .......... .......... .......... .......... .......... 42%  345M 2s
  2400K .......... .......... .......... .......... .......... 43% 30.2M 1s
  2450K .......... .......... .......... .......... .......... 44%  216M 1s
  2500K .......... .......... .......... .......... .......... 45% 4.64M 1s
  2550K .......... .......... .......... .......... .......... 46%  128M 1s
  2600K .......... .......... .......... .......... .......... 47%  620M 1s
  2650K .......... .......... .......... .......... .......... 47%  135M 1s
  2700K .......... .......... .......... .......... .......... 48%  186M 1s
  2750K .......... .......... .......... .......... .......... 49% 96.0M 1s
  2800K .......... .......... .......... .......... .......... 50%  628M 1s
  2850K .......... .......... .......... .......... .......... 51%  158M 1s
  2900K .......... .......... .......... .......... .......... 52%  256M 1s
  2950K .......... .......... .......... .......... .......... 53%  553M 1s
  3000K .......... .......... .......... .......... .......... 54%  247M 1s
  3050K .......... .......... .......... .......... .......... 55%  190M 1s
  3100K .......... .......... .......... .......... .......... 55%  311M 1s
  3150K .......... .......... .......... .......... .......... 56%  488M 1s
  3200K .......... .......... .......... .......... .......... 57%  614M 1s
  3250K .......... .......... .......... .......... .......... 58%  104M 1s
  3300K .......... .......... .......... .......... .......... 59%  303M 1s
  3350K .......... .......... .......... .......... .......... 60%  103M 1s
  3400K .......... .......... .......... .......... .......... 61%  112M 1s
  3450K .......... .......... .......... .......... .......... 62% 4.85M 1s
  3500K .......... .......... .......... .......... .......... 63%  208M 1s
  3550K .......... .......... .......... .......... .......... 63%  290M 1s
  3600K .......... .......... .......... .......... .......... 64%  343M 1s
  3650K .......... .......... .......... .......... .......... 65%  137M 1s
  3700K .......... .......... .......... .......... .......... 66%  349M 1s
  3750K .......... .......... .......... .......... .......... 67%  201M 1s
  3800K .......... .......... .......... .......... .......... 68%  212M 1s
  3850K .......... .......... .......... .......... .......... 69%  295M 1s
  3900K .......... .......... .......... .......... .......... 70%  483M 1s
  3950K .......... .......... .......... .......... .......... 71%  396M 1s
  4000K .......... .......... .......... .......... .......... 71%  274M 1s
  4050K .......... .......... .......... .......... .......... 72%  169M 1s
  4100K .......... .......... .......... .......... .......... 73%  580M 0s
  4150K .......... .......... .......... .......... .......... 74%  198M 0s
  4200K .......... .......... .......... .......... .......... 75%  367M 0s
  4250K .......... .......... .......... .......... .......... 76%  593M 0s
  4300K .......... .......... .......... .......... .......... 77%  201M 0s
  4350K .......... .......... .......... .......... .......... 78%  298M 0s
  4400K .......... .......... .......... .......... .......... 79%  505M 0s
  4450K .......... .......... .......... .......... .......... 79%  336M 0s
  4500K .......... .......... .......... .......... .......... 80%  245M 0s
  4550K .......... .......... .......... .......... .......... 81%  285M 0s
  4600K .......... .......... .......... .......... .......... 82%  283M 0s
  4650K .......... .......... .......... .......... .......... 83%  280M 0s
  4700K .......... .......... .......... .......... .......... 84%  435M 0s
  4750K .......... .......... .......... .......... .......... 85%  246M 0s
  4800K .......... .......... .......... .......... .......... 86%  306M 0s
  4850K .......... .......... .......... .......... .......... 87%  206M 0s
  4900K .......... .......... .......... .......... .......... 87%  273M 0s
  4950K .......... .......... .......... .......... .......... 88% 3.01M 0s
  5000K .......... .......... .......... .......... .......... 89%  186M 0s
  5050K .......... .......... .......... .......... .......... 90% 1.12G 0s
  5100K .......... .......... .......... .......... .......... 91% 1.53G 0s
  5150K .......... .......... .......... .......... .......... 92% 1.55G 0s
  5200K .......... .......... .......... .......... .......... 93% 1.07G 0s
  5250K .......... .......... .......... .......... .......... 94% 1.76G 0s
  5300K .......... .......... .......... .......... .......... 95% 1.04G 0s
  5350K .......... .......... .......... .......... .......... 95% 2.08G 0s
  5400K .......... .......... .......... .......... .......... 96% 1.58G 0s
  5450K .......... .......... .......... .......... .......... 97% 1.24G 0s
  5500K .......... .......... .......... .......... .......... 98% 1.90G 0s
  5550K .......... .......... .......... .......... .......... 99% 2.38G 0s
  5600K .......... .......... .......... .                    100% 2.43G=1.5s

2020-03-02 03:27:18 (30.0 Mb/s) - ‘/dev/null’ saved [5766625/5766625]

