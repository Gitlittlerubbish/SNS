--2020-03-02 03:24:02--  http://www.mined.gob.sv/sexualidad/Media.pdf
Resolving www.mined.gob.sv (www.mined.gob.sv)... 168.243.116.34
Connecting to www.mined.gob.sv (www.mined.gob.sv)|168.243.116.34|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 4552975 (4.3M) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  1% 1.31M 28s
    50K .......... .......... .......... .......... ..........  2% 2.63M 20s
   100K .......... .......... .......... .......... ..........  3% 86.5M 14s
   150K .......... .......... .......... .......... ..........  4%  160M 10s
   200K .......... .......... .......... .......... ..........  5% 2.71M 11s
   250K .......... .......... .......... .......... ..........  6% 56.1M 9s
   300K .......... .......... .......... .......... ..........  7% 2.73M 9s
   350K .......... .......... .......... .......... ..........  8%  156M 8s
   400K .......... .......... .......... .......... .......... 10%  338M 7s
   450K .......... .......... .......... .......... .......... 11%  309M 6s
   500K .......... .......... .......... .......... .......... 12%  115M 6s
   550K .......... .......... .......... .......... .......... 13% 2.74M 6s
   600K .......... .......... .......... .......... .......... 14%  117M 6s
   650K .......... .......... .......... .......... .......... 15% 80.5M 5s
   700K .......... .......... .......... .......... .......... 16%  647M 5s
   750K .......... .......... .......... .......... .......... 17% 2.85M 5s
   800K .......... .......... .......... .......... .......... 19%  134M 5s
   850K .......... .......... .......... .......... .......... 20% 1.09G 4s
   900K .......... .......... .......... .......... .......... 21%  153M 4s
   950K .......... .......... .......... .......... .......... 22%  188M 4s
  1000K .......... .......... .......... .......... .......... 23%  267M 4s
  1050K .......... .......... .......... .......... .......... 24%  128M 3s
  1100K .......... .......... .......... .......... .......... 25%  131M 3s
  1150K .......... .......... .......... .......... .......... 26% 4.01M 3s
  1200K .......... .......... .......... .......... .......... 28% 9.91M 3s
  1250K .......... .......... .......... .......... .......... 29%  191M 3s
  1300K .......... .......... .......... .......... .......... 30%  155M 3s
  1350K .......... .......... .......... .......... .......... 31%  250M 3s
  1400K .......... .......... .......... .......... .......... 32%  126M 3s
  1450K .......... .......... .......... .......... .......... 33%  340M 2s
  1500K .......... .......... .......... .......... .......... 34%  246M 2s
  1550K .......... .......... .......... .......... .......... 35%  221M 2s
  1600K .......... .......... .......... .......... .......... 37%  196M 2s
  1650K .......... .......... .......... .......... .......... 38% 4.08M 2s
  1700K .......... .......... .......... .......... .......... 39% 9.75M 2s
  1750K .......... .......... .......... .......... .......... 40%  121M 2s
  1800K .......... .......... .......... .......... .......... 41%  355M 2s
  1850K .......... .......... .......... .......... .......... 42%  290M 2s
  1900K .......... .......... .......... .......... .......... 43%  241M 2s
  1950K .......... .......... .......... .......... .......... 44%  352M 2s
  2000K .......... .......... .......... .......... .......... 46%  235M 2s
  2050K .......... .......... .......... .......... .......... 47%  332M 2s
  2100K .......... .......... .......... .......... .......... 48%  328M 2s
  2150K .......... .......... .......... .......... .......... 49%  225M 1s
  2200K .......... .......... .......... .......... .......... 50%  484M 1s
  2250K .......... .......... .......... .......... .......... 51%  540M 1s
  2300K .......... .......... .......... .......... .......... 52%  343M 1s
  2350K .......... .......... .......... .......... .......... 53%  234M 1s
  2400K .......... .......... .......... .......... .......... 55%  335M 1s
  2450K .......... .......... .......... .......... .......... 56% 4.45M 1s
  2500K .......... .......... .......... .......... .......... 57% 9.34M 1s
  2550K .......... .......... .......... .......... .......... 58%  130M 1s
  2600K .......... .......... .......... .......... .......... 59%  623M 1s
  2650K .......... .......... .......... .......... .......... 60% 85.8M 1s
  2700K .......... .......... .......... .......... .......... 61%  716M 1s
  2750K .......... .......... .......... .......... .......... 62%  387M 1s
  2800K .......... .......... .......... .......... .......... 64%  150M 1s
  2850K .......... .......... .......... .......... .......... 65% 36.2M 1s
  2900K .......... .......... .......... .......... .......... 66%  112M 1s
  2950K .......... .......... .......... .......... .......... 67%  317M 1s
  3000K .......... .......... .......... .......... .......... 68% 65.6M 1s
  3050K .......... .......... .......... .......... .......... 69% 97.3M 1s
  3100K .......... .......... .......... .......... .......... 70%  147M 1s
  3150K .......... .......... .......... .......... .......... 71%  197M 1s
  3200K .......... .......... .......... .......... .......... 73%  166M 1s
  3250K .......... .......... .......... .......... .......... 74% 8.65M 1s
  3300K .......... .......... .......... .......... .......... 75% 33.9M 1s
  3350K .......... .......... .......... .......... .......... 76%  153M 1s
  3400K .......... .......... .......... .......... .......... 77%  104M 0s
  3450K .......... .......... .......... .......... .......... 78% 87.6M 0s
  3500K .......... .......... .......... .......... .......... 79% 7.42M 0s
  3550K .......... .......... .......... .......... .......... 80% 48.7M 0s
  3600K .......... .......... .......... .......... .......... 82%  118M 0s
  3650K .......... .......... .......... .......... .......... 83%  495M 0s
  3700K .......... .......... .......... .......... .......... 84% 69.0M 0s
  3750K .......... .......... .......... .......... .......... 85%  271M 0s
  3800K .......... .......... .......... .......... .......... 86%  169M 0s
  3850K .......... .......... .......... .......... .......... 87%  661M 0s
  3900K .......... .......... .......... .......... .......... 88%  358M 0s
  3950K .......... .......... .......... .......... .......... 89%  222M 0s
  4000K .......... .......... .......... .......... .......... 91%  389M 0s
  4050K .......... .......... .......... .......... .......... 92%  306M 0s
  4100K .......... .......... .......... .......... .......... 93%  121M 0s
  4150K .......... .......... .......... .......... .......... 94%  366M 0s
  4200K .......... .......... .......... .......... .......... 95%  172M 0s
  4250K .......... .......... .......... .......... .......... 96%  111M 0s
  4300K .......... .......... .......... .......... .......... 97%  450M 0s
  4350K .......... .......... .......... .......... .......... 98%  209M 0s
  4400K .......... .......... .......... .......... ......    100% 10.0M=1.8s

2020-03-02 03:24:05 (20.0 Mb/s) - ‘/dev/null’ saved [4552975/4552975]

