--2020-02-25 22:14:18--  http://www.censos.gob.sv/cpv/descargas/CPV_Proyeccion_Resultados.pdf%0D
Resolving www.censos.gob.sv (www.censos.gob.sv)... 200.89.85.145
Connecting to www.censos.gob.sv (www.censos.gob.sv)|200.89.85.145|:80... connected.
HTTP request sent, awaiting response... 400 Bad Request
2020-02-25 22:14:19 ERROR 400: Bad Request.

--2020-02-25 22:14:39--  http://www.censos.gob.sv/cpv/descargas/CPV_Proyeccion_Resultados.pdf%0D
Resolving www.censos.gob.sv (www.censos.gob.sv)... 200.89.85.145
Connecting to www.censos.gob.sv (www.censos.gob.sv)|200.89.85.145|:80... connected.
HTTP request sent, awaiting response... 400 Bad Request
2020-02-25 22:14:39 ERROR 400: Bad Request.

