--2020-02-25 22:12:41--  http://www.ufg.edu.sv/doc/FT-EBSCOhost.pdf%0D
Resolving www.ufg.edu.sv (www.ufg.edu.sv)... 200.124.138.25
Connecting to www.ufg.edu.sv (www.ufg.edu.sv)|200.124.138.25|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:12:43 ERROR 404: Not Found.

--2020-02-25 22:13:22--  http://www.ufg.edu.sv/doc/FT-EBSCOhost.pdf%0D
Resolving www.ufg.edu.sv (www.ufg.edu.sv)... 200.124.138.25
Connecting to www.ufg.edu.sv (www.ufg.edu.sv)|200.124.138.25|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:22 ERROR 404: Not Found.

