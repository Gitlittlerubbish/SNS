--2020-03-02 03:24:07--  http://richmond.com.sv/ss/SSpathwaytoscience_g.pdf
Resolving richmond.com.sv (richmond.com.sv)... 34.225.172.62, 34.238.101.91
Connecting to richmond.com.sv (richmond.com.sv)|34.225.172.62|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 429661 (420K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 11% 2.38M 1s
    50K .......... .......... .......... .......... .......... 23% 4.80M 1s
   100K .......... .......... .......... .......... .......... 35%  134M 0s
   150K .......... .......... .......... .......... .......... 47% 93.8M 0s
   200K .......... .......... .......... .......... .......... 59% 5.03M 0s
   250K .......... .......... .......... .......... .......... 71% 99.0M 0s
   300K .......... .......... .......... .......... .......... 83% 5.13M 0s
   350K .......... .......... .......... .......... .......... 95%  145M 0s
   400K .......... .........                                  100% 1.71G=0.4s

2020-03-02 03:24:07 (7.94 Mb/s) - ‘/dev/null’ saved [429661/429661]

