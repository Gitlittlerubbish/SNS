--2020-02-25 22:12:55--  https://www.cortedecuentas.gob.sv/genero/PROTOCOLO.pdf%0D
Resolving www.cortedecuentas.gob.sv (www.cortedecuentas.gob.sv)... 190.5.130.194
Connecting to www.cortedecuentas.gob.sv (www.cortedecuentas.gob.sv)|190.5.130.194|:443... connected.
HTTP request sent, awaiting response... 500 Internal Server Error
2020-02-25 22:12:56 ERROR 500: Internal Server Error.

--2020-02-25 22:12:56--  https://www.cortedecuentas.gob.sv/images/ccrevista.pdf%0D
Resolving www.cortedecuentas.gob.sv (www.cortedecuentas.gob.sv)... 190.5.130.194
Connecting to www.cortedecuentas.gob.sv (www.cortedecuentas.gob.sv)|190.5.130.194|:443... connected.
HTTP request sent, awaiting response... 500 Internal Server Error
2020-02-25 22:12:56 ERROR 500: Internal Server Error.

--2020-02-25 22:13:31--  https://www.cortedecuentas.gob.sv/genero/PROTOCOLO.pdf%0D
Resolving www.cortedecuentas.gob.sv (www.cortedecuentas.gob.sv)... 190.5.130.194
Connecting to www.cortedecuentas.gob.sv (www.cortedecuentas.gob.sv)|190.5.130.194|:443... connected.
HTTP request sent, awaiting response... 500 Internal Server Error
2020-02-25 22:13:31 ERROR 500: Internal Server Error.

--2020-02-25 22:13:31--  https://www.cortedecuentas.gob.sv/images/ccrevista.pdf%0D
Resolving www.cortedecuentas.gob.sv (www.cortedecuentas.gob.sv)... 190.5.130.194
Connecting to www.cortedecuentas.gob.sv (www.cortedecuentas.gob.sv)|190.5.130.194|:443... connected.
HTTP request sent, awaiting response... 500 Internal Server Error
2020-02-25 22:13:32 ERROR 500: Internal Server Error.

