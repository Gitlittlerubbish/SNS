--2020-02-25 22:13:01--  https://thyssenkrupp.com.sv/noticia/download/763/%0D
Resolving thyssenkrupp.com.sv (thyssenkrupp.com.sv)... 186.202.143.17
Connecting to thyssenkrupp.com.sv (thyssenkrupp.com.sv)|186.202.143.17|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: 1282642 (1.2M) [application/download]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  3%  536K 18s
    50K .......... .......... .......... .......... ..........  7%  804K 15s
   100K .......... .......... .......... .......... .......... 11% 11.0M 10s
   150K .......... .......... .......... .......... .......... 15% 1.59M 8s
   200K .......... .......... .......... .......... .......... 19% 1.91M 7s
   250K .......... .......... .......... .......... .......... 23% 1.61M 6s
   300K .......... .......... .......... .......... .......... 27% 1.61M 6s
   350K .......... .......... .......... .......... .......... 31%  431K 7s
   400K .......... .......... .......... .......... .......... 35%  537K 7s
   450K .......... .......... .......... .......... .......... 39%  805K 7s
   500K .......... .......... .......... .......... .......... 43%  403K 7s
   550K .......... .......... .......... .......... .......... 47%  179K 9s
   600K .......... .......... .......... .......... .......... 51%  403K 8s
   650K .......... .......... .......... .......... .......... 55%  537K 8s
   700K .......... .......... .......... .......... .......... 59%  537K 7s
   750K .......... .......... .......... .......... .......... 63%  805K 6s
   800K .......... .......... .......... .......... .......... 67%  804K 5s
   850K .......... .......... .......... .......... .......... 71%  804K 5s
   900K .......... .......... .......... .......... .......... 75% 1.61M 4s
   950K .......... .......... .......... .......... .......... 79%  805K 3s
  1000K .......... .......... .......... .......... .......... 83%  322K 3s
  1050K .......... .......... .......... .......... .......... 87%  403K 2s
  1100K .......... .......... .......... .......... .......... 91%  805K 1s
  1150K .......... .......... .......... .......... .......... 95%  537K 1s
  1200K .......... .......... .......... .......... .......... 99% 1.61M 0s
  1250K ..                                                    100% 42272G=16s

2020-02-25 22:13:19 (623 Kb/s) - ‘/dev/null’ saved [1282642/1282642]

--2020-02-25 22:13:19--  https://thyssenkrupp.com.sv/noticia/download/763/%0D
Resolving thyssenkrupp.com.sv (thyssenkrupp.com.sv)... 186.202.143.17
Connecting to thyssenkrupp.com.sv (thyssenkrupp.com.sv)|186.202.143.17|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: 1282642 (1.2M) [application/download]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  3%  532K 19s
    50K .......... .......... .......... .......... ..........  7% 1.38M 12s
   100K .......... .......... .......... .......... .......... 11% 1.90M 9s
   150K .......... .......... .......... .......... .......... 15% 1.60M 8s
   200K .......... .......... .......... .......... .......... 19% 1.60M 7s
   250K .......... .......... .......... .......... .......... 23%  399K 9s
   300K .......... .......... .......... .......... .......... 27%  798K 9s
   350K .......... .......... .......... .......... .......... 31% 1.38M 8s
   400K .......... .......... .......... .......... .......... 35%  867K 7s
   450K .......... .......... .......... .......... .......... 39% 1.38M 7s
   500K .......... .......... .......... .......... .......... 43% 1.60M 6s
   550K .......... .......... .......... .......... .......... 47% 1.60M 5s
   600K .......... .......... .......... .......... .......... 51%  233K 6s
   650K .......... .......... .......... .......... .......... 55%  743K 6s
   700K .......... .......... .......... .......... .......... 59%  560K 5s
   750K .......... .......... .......... .......... .......... 63% 1.59M 5s
   800K .......... .......... .......... .......... .......... 67%  798K 4s
   850K .......... .......... .......... .......... .......... 71% 1.60M 4s
   900K .......... .......... .......... .......... .......... 75%  798K 3s
   950K .......... .......... .......... .......... .......... 79%  399K 3s
  1000K .......... .......... .......... .......... .......... 83%  532K 2s
  1050K .......... .......... .......... .......... .......... 87%  532K 2s
  1100K .......... .......... .......... .......... .......... 91%  798K 1s
  1150K .......... .......... .......... .......... .......... 95%  798K 1s
  1200K .......... .......... .......... .......... .......... 99% 1.60M 0s
  1250K ..                                                    100% 42272G=13s

2020-02-25 22:13:34 (769 Kb/s) - ‘/dev/null’ saved [1282642/1282642]

--2020-02-25 22:13:35--  https://thyssenkrupp.com.sv/noticia/download/763/%0D
Resolving thyssenkrupp.com.sv (thyssenkrupp.com.sv)... 186.202.143.17
Connecting to thyssenkrupp.com.sv (thyssenkrupp.com.sv)|186.202.143.17|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: 1282642 (1.2M) [application/download]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  3%  532K 19s
    50K .......... .......... .......... .......... ..........  7%  799K 15s
   100K .......... .......... .......... .......... .......... 11%  798K 13s
   150K .......... .......... .......... .......... .......... 15%  798K 12s
   200K .......... .......... .......... .......... .......... 19%  266K 15s
   250K .......... .......... .......... .......... .......... 23%  532K 15s
   300K .......... .......... .......... .......... .......... 27%  532K 14s
   350K .......... .......... .......... .......... .......... 31% 1.60M 12s
   400K .......... .......... .......... .......... .......... 35%  799K 11s
   450K .......... .......... .......... .......... .......... 39%  266K 12s
   500K .......... .......... .......... .......... .......... 43%  532K 11s
   550K .......... .......... .......... .......... .......... 47%  532K 10s
   600K .......... .......... .......... .......... .......... 51%  798K 9s
   650K .......... .......... .......... .......... .......... 55%  798K 8s
   700K .......... .......... .......... .......... .......... 59%  266K 8s
   750K .......... .......... .......... .......... .......... 63%  798K 7s
   800K .......... .......... .......... .......... .......... 67%  532K 6s
   850K .......... .......... .......... .......... .......... 71%  798K 5s
   900K .......... .......... .......... .......... .......... 75%  228K 5s
   950K .......... .......... .......... .......... .......... 79%  399K 4s
  1000K .......... .......... .......... .......... .......... 83%  532K 3s
  1050K .......... .......... .......... .......... .......... 87%  532K 2s
  1100K .......... .......... .......... .......... .......... 91%  798K 2s
  1150K .......... .......... .......... .......... .......... 95% 1.60M 1s
  1200K .......... .......... .......... .......... .......... 99%  797K 0s
  1250K ..                                                    100% 42272G=19s

2020-02-25 22:13:55 (533 Kb/s) - ‘/dev/null’ saved [1282642/1282642]

--2020-02-25 22:13:55--  https://thyssenkrupp.com.sv/noticia/download/763/%0D
Resolving thyssenkrupp.com.sv (thyssenkrupp.com.sv)... 186.202.143.17
Connecting to thyssenkrupp.com.sv (thyssenkrupp.com.sv)|186.202.143.17|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: 1282642 (1.2M) [application/download]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  3%  543K 18s
    50K .......... .......... .......... .......... ..........  7%  814K 14s
   100K .......... .......... .......... .......... .......... 11%  815K 13s
   150K .......... .......... .......... .......... .......... 15%  815K 12s
   200K .......... .......... .......... .......... .......... 19% 1.63M 10s
   250K .......... .......... .......... .......... .......... 23%  814K 10s
   300K .......... .......... .......... .......... .......... 27% 1.63M 8s
   350K .......... .......... .......... .......... .......... 31%  815K 8s
   400K .......... .......... .......... .......... .......... 35%  272K 9s
   450K .......... .......... .......... .......... .......... 39%  543K 9s
   500K .......... .......... .......... .......... .......... 43%  814K 8s
   550K .......... .......... .......... .......... .......... 47%  815K 8s
   600K .......... .......... .......... .......... .......... 51%  814K 7s
   650K .......... .......... .......... .......... .......... 55% 1.63M 6s
   700K .......... .......... .......... .......... .......... 59%  815K 6s
   750K .......... .......... .......... .......... .......... 63%  909K 5s
   800K .......... .......... .......... .......... .......... 67% 1.35M 4s
   850K .......... .......... .......... .......... .......... 71% 1.63M 4s
   900K .......... .......... .......... .......... .......... 75% 1.63M 3s
   950K .......... .......... .......... .......... .......... 79%  815K 3s
  1000K .......... .......... .......... .......... .......... 83% 1.63M 2s
  1050K .......... .......... .......... .......... .......... 87% 1.63M 1s
  1100K .......... .......... .......... .......... .......... 91% 1.63M 1s
  1150K .......... .......... .......... .......... .......... 95% 1.63M 0s
  1200K .......... .......... .......... .......... .......... 99% 1.63M 0s
  1250K ..                                                    100% 42272G=11s

2020-02-25 22:14:08 (907 Kb/s) - ‘/dev/null’ saved [1282642/1282642]

