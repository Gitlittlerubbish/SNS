--2020-02-25 22:13:35--  http://www.cultura.gob.sv/wp-content/uploads/2016/08/Revista_ARS_10.pdf%0D
Resolving www.cultura.gob.sv (www.cultura.gob.sv)... 190.120.4.18
Connecting to www.cultura.gob.sv (www.cultura.gob.sv)|190.120.4.18|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:39 ERROR 404: Not Found.

--2020-02-25 22:14:08--  http://www.cultura.gob.sv/wp-content/uploads/2016/08/Revista_ARS_10.pdf%0D
Resolving www.cultura.gob.sv (www.cultura.gob.sv)... 190.120.4.18
Connecting to www.cultura.gob.sv (www.cultura.gob.sv)|190.120.4.18|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:09 ERROR 404: Not Found.

