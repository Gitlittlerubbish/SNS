--2020-02-25 22:13:42--  http://puntosdeventa.com.sv/manuales/47/DS000003_1515L.pdf%0D
Resolving puntosdeventa.com.sv (puntosdeventa.com.sv)... 67.227.226.242
Connecting to puntosdeventa.com.sv (puntosdeventa.com.sv)|67.227.226.242|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:42 ERROR 404: Not Found.

--2020-02-25 22:14:11--  http://puntosdeventa.com.sv/manuales/47/DS000003_1515L.pdf%0D
Resolving puntosdeventa.com.sv (puntosdeventa.com.sv)... 67.227.226.242
Connecting to puntosdeventa.com.sv (puntosdeventa.com.sv)|67.227.226.242|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:11 ERROR 404: Not Found.

