--2020-02-25 22:12:52--  http://www.fiaes.org.sv/library/desarrolloterritorialysostenibilidadambiental.pdf%0D
Resolving www.fiaes.org.sv (www.fiaes.org.sv)... 95.216.100.230
Connecting to www.fiaes.org.sv (www.fiaes.org.sv)|95.216.100.230|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: https://www.fiaes.org.sv/library/desarrolloterritorialysostenibilidadambiental.pdf%0d [following]
--2020-02-25 22:12:52--  https://www.fiaes.org.sv/library/desarrolloterritorialysostenibilidadambiental.pdf%0d
Connecting to www.fiaes.org.sv (www.fiaes.org.sv)|95.216.100.230|:443... connected.
HTTP request sent, awaiting response... 404 NOT FOUND
2020-02-25 22:12:52 ERROR 404: NOT FOUND.

--2020-02-25 22:13:28--  http://www.fiaes.org.sv/library/desarrolloterritorialysostenibilidadambiental.pdf%0D
Resolving www.fiaes.org.sv (www.fiaes.org.sv)... 95.216.100.230
Connecting to www.fiaes.org.sv (www.fiaes.org.sv)|95.216.100.230|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: https://www.fiaes.org.sv/library/desarrolloterritorialysostenibilidadambiental.pdf%0d [following]
--2020-02-25 22:13:28--  https://www.fiaes.org.sv/library/desarrolloterritorialysostenibilidadambiental.pdf%0d
Connecting to www.fiaes.org.sv (www.fiaes.org.sv)|95.216.100.230|:443... connected.
HTTP request sent, awaiting response... 404 NOT FOUND
2020-02-25 22:13:28 ERROR 404: NOT FOUND.

