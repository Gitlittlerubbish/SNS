--2020-02-25 22:12:50--  http://www.fundar.org.sv/referencias/pipilpots.pdf%0D
Resolving www.fundar.org.sv (www.fundar.org.sv)... 190.120.10.123
Connecting to www.fundar.org.sv (www.fundar.org.sv)|190.120.10.123|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:12:50 ERROR 404: Not Found.

--2020-02-25 22:13:27--  http://www.fundar.org.sv/referencias/pipilpots.pdf%0D
Resolving www.fundar.org.sv (www.fundar.org.sv)... 190.120.10.123
Connecting to www.fundar.org.sv (www.fundar.org.sv)|190.120.10.123|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:27 ERROR 404: Not Found.

