--2020-03-02 03:23:47--  http://www.marn.gob.sv/inema2017.pdf
Resolving www.marn.gob.sv (www.marn.gob.sv)... 104.210.5.96
Connecting to www.marn.gob.sv (www.marn.gob.sv)|104.210.5.96|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 36499294 (35M) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  0% 2.48M 1m58s
    50K .......... .......... .......... .......... ..........  0% 4.95M 88s
   100K .......... .......... .......... .......... ..........  0%  115M 60s
   150K .......... .......... .......... .......... ..........  0%  159M 45s
   200K .......... .......... .......... .......... ..........  0% 4.97M 48s
   250K .......... .......... .......... .......... ..........  0%  185M 40s
   300K .......... .......... .......... .......... ..........  0% 5.32M 42s
   350K .......... .......... .......... .......... ..........  1%  235M 37s
   400K .......... .......... .......... .......... ..........  1%  422M 33s
   450K .......... .......... .......... .......... ..........  1%  110M 30s
   500K .......... .......... .......... .......... ..........  1%  229M 27s
   550K .......... .......... .......... .......... ..........  1% 5.32M 29s
   600K .......... .......... .......... .......... ..........  1%  114M 27s
   650K .......... .......... .......... .......... ..........  1%  237M 25s
   700K .......... .......... .......... .......... ..........  2%  101M 24s
   750K .......... .......... .......... .......... ..........  2%  464M 22s
   800K .......... .......... .......... .......... ..........  2% 5.57M 24s
   850K .......... .......... .......... .......... ..........  2%  268M 23s
   900K .......... .......... .......... .......... ..........  2%  342M 21s
   950K .......... .......... .......... .......... ..........  2%  369M 20s
  1000K .......... .......... .......... .......... ..........  2%  229M 19s
  1050K .......... .......... .......... .......... ..........  3%  408M 19s
  1100K .......... .......... .......... .......... ..........  3%  109M 18s
  1150K .......... .......... .......... .......... ..........  3%  421M 17s
  1200K .......... .......... .......... .......... ..........  3% 5.30M 19s
  1250K .......... .......... .......... .......... ..........  3%  136M 18s
  1300K .......... .......... .......... .......... ..........  3%  340M 17s
  1350K .......... .......... .......... .......... ..........  3%  138M 17s
  1400K .......... .......... .......... .......... ..........  4%  720M 16s
  1450K .......... .......... .......... .......... ..........  4%  328M 16s
  1500K .......... .......... .......... .......... ..........  4%  314M 15s
  1550K .......... .......... .......... .......... ..........  4%  231M 15s
  1600K .......... .......... .......... .......... ..........  4%  226M 14s
  1650K .......... .......... .......... .......... ..........  4% 6.07M 15s
  1700K .......... .......... .......... .......... ..........  4%  159M 15s
  1750K .......... .......... .......... .......... ..........  5%  320M 14s
  1800K .......... .......... .......... .......... ..........  5%  237M 14s
  1850K .......... .......... .......... .......... ..........  5%  292M 14s
  1900K .......... .......... .......... .......... ..........  5%  253M 13s
  1950K .......... .......... .......... .......... ..........  5%  492M 13s
  2000K .......... .......... .......... .......... ..........  5%  346M 13s
  2050K .......... .......... .......... .......... ..........  5%  225M 12s
  2100K .......... .......... .......... .......... ..........  6%  380M 12s
  2150K .......... .......... .......... .......... ..........  6%  212M 12s
  2200K .......... .......... .......... .......... ..........  6%  223M 11s
  2250K .......... .......... .......... .......... ..........  6%  265M 11s
  2300K .......... .......... .......... .......... ..........  6%  735M 11s
  2350K .......... .......... .......... .......... ..........  6%  281M 11s
  2400K .......... .......... .......... .......... ..........  6%  171M 11s
  2450K .......... .......... .......... .......... ..........  7%  163M 10s
  2500K .......... .......... .......... .......... ..........  7% 6.92M 11s
  2550K .......... .......... .......... .......... ..........  7%  103M 11s
  2600K .......... .......... .......... .......... ..........  7% 87.7M 11s
  2650K .......... .......... .......... .......... ..........  7%  201M 10s
  2700K .......... .......... .......... .......... ..........  7%  423M 10s
  2750K .......... .......... .......... .......... ..........  7%  283M 10s
  2800K .......... .......... .......... .......... ..........  7%  272M 10s
  2850K .......... .......... .......... .......... ..........  8%  155M 10s
  2900K .......... .......... .......... .......... ..........  8%  412M 10s
  2950K .......... .......... .......... .......... ..........  8%  187M 9s
  3000K .......... .......... .......... .......... ..........  8%  389M 9s
  3050K .......... .......... .......... .......... ..........  8%  345M 9s
  3100K .......... .......... .......... .......... ..........  8%  196M 9s
  3150K .......... .......... .......... .......... ..........  8%  344M 9s
  3200K .......... .......... .......... .......... ..........  9%  241M 9s
  3250K .......... .......... .......... .......... ..........  9%  146M 9s
  3300K .......... .......... .......... .......... ..........  9%  353M 8s
  3350K .......... .......... .......... .......... ..........  9% 8.07M 9s
  3400K .......... .......... .......... .......... ..........  9%  343M 9s
  3450K .......... .......... .......... .......... ..........  9%  191M 8s
  3500K .......... .......... .......... .......... ..........  9%  481M 8s
  3550K .......... .......... .......... .......... .......... 10%  438M 8s
  3600K .......... .......... .......... .......... .......... 10%  214M 8s
  3650K .......... .......... .......... .......... .......... 10%  350M 8s
  3700K .......... .......... .......... .......... .......... 10%  223M 8s
  3750K .......... .......... .......... .......... .......... 10%  332M 8s
  3800K .......... .......... .......... .......... .......... 10%  584M 8s
  3850K .......... .......... .......... .......... .......... 10% 86.7M 8s
  3900K .......... .......... .......... .......... .......... 11%  226M 8s
  3950K .......... .......... .......... .......... .......... 11%  198M 7s
  4000K .......... .......... .......... .......... .......... 11%  453M 7s
  4050K .......... .......... .......... .......... .......... 11% 2.25M 9s
  4100K .......... .......... .......... .......... .......... 11% 1.91G 9s
  4150K .......... .......... .......... .......... .......... 11%  256M 8s
  4200K .......... .......... .......... .......... .......... 11%  175M 8s
  4250K .......... .......... .......... .......... .......... 12% 1.78G 8s
  4300K .......... .......... .......... .......... .......... 12% 1.02G 8s
  4350K .......... .......... .......... .......... .......... 12% 91.7M 8s
  4400K .......... .......... .......... .......... .......... 12%  163M 8s
  4450K .......... .......... .......... .......... .......... 12% 2.13G 8s
  4500K .......... .......... .......... .......... .......... 12% 1.46G 8s
  4550K .......... .......... .......... .......... .......... 12% 2.16G 8s
  4600K .......... .......... .......... .......... .......... 13% 2.51G 8s
  4650K .......... .......... .......... .......... .......... 13% 2.18G 7s
  4700K .......... .......... .......... .......... .......... 13% 2.53G 7s
  4750K .......... .......... .......... .......... .......... 13% 2.54G 7s
  4800K .......... .......... .......... .......... .......... 13% 2.53G 7s
  4850K .......... .......... .......... .......... .......... 13% 2.18G 7s
  4900K .......... .......... .......... .......... .......... 13% 2.53G 7s
  4950K .......... .......... .......... .......... .......... 14% 2.40G 7s
  5000K .......... .......... .......... .......... .......... 14% 2.28G 7s
  5050K .......... .......... .......... .......... .......... 14% 1.93G 7s
  5100K .......... .......... .......... .......... .......... 14% 3.15G 7s
  5150K .......... .......... .......... .......... .......... 14% 2.54G 7s
  5200K .......... .......... .......... .......... .......... 14% 3.30G 7s
  5250K .......... .......... .......... .......... .......... 14% 2.53G 7s
  5300K .......... .......... .......... .......... .......... 15% 3.18G 6s
  5350K .......... .......... .......... .......... .......... 15% 3.25G 6s
  5400K .......... .......... .......... .......... .......... 15%  119M 6s
  5450K .......... .......... .......... .......... .......... 15%  189M 6s
  5500K .......... .......... .......... .......... .......... 15%  104M 6s
  5550K .......... .......... .......... .......... .......... 15%  352M 6s
  5600K .......... .......... .......... .......... .......... 15%  120M 6s
  5650K .......... .......... .......... .......... .......... 15% 12.5M 6s
  5700K .......... .......... .......... .......... .......... 16%  265M 6s
  5750K .......... .......... .......... .......... .......... 16% 19.7M 6s
  5800K .......... .......... .......... .......... .......... 16%  270M 6s
  5850K .......... .......... .......... .......... .......... 16%  184M 6s
  5900K .......... .......... .......... .......... .......... 16%  261M 6s
  5950K .......... .......... .......... .......... .......... 16%  409M 6s
  6000K .......... .......... .......... .......... .......... 16%  151M 6s
  6050K .......... .......... .......... .......... .......... 17% 1.17G 6s
  6100K .......... .......... .......... .......... .......... 17%  103M 6s
  6150K .......... .......... .......... .......... .......... 17%  379M 6s
  6200K .......... .......... .......... .......... .......... 17%  481M 6s
  6250K .......... .......... .......... .......... .......... 17%  224M 6s
  6300K .......... .......... .......... .......... .......... 17%  273M 6s
  6350K .......... .......... .......... .......... .......... 17%  407M 6s
  6400K .......... .......... .......... .......... .......... 18%  406M 6s
  6450K .......... .......... .......... .......... .......... 18%  150M 6s
  6500K .......... .......... .......... .......... .......... 18%  212M 5s
  6550K .......... .......... .......... .......... .......... 18%  300M 5s
  6600K .......... .......... .......... .......... .......... 18%  168M 5s
  6650K .......... .......... .......... .......... .......... 18% 12.7M 5s
  6700K .......... .......... .......... .......... .......... 18%  175M 5s
  6750K .......... .......... .......... .......... .......... 19%  457M 5s
  6800K .......... .......... .......... .......... .......... 19%  481M 5s
  6850K .......... .......... .......... .......... .......... 19%  192M 5s
  6900K .......... .......... .......... .......... .......... 19%  451M 5s
  6950K .......... .......... .......... .......... .......... 19%  165M 5s
  7000K .......... .......... .......... .......... .......... 19% 67.0M 5s
  7050K .......... .......... .......... .......... .......... 19% 1.55M 6s
  7100K .......... .......... .......... .......... .......... 20% 1.36G 6s
  7150K .......... .......... .......... .......... .......... 20% 1.65G 6s
  7200K .......... .......... .......... .......... .......... 20% 1.83G 6s
  7250K .......... .......... .......... .......... .......... 20% 1.89G 6s
  7300K .......... .......... .......... .......... .......... 20% 1.77G 6s
  7350K .......... .......... .......... .......... .......... 20% 1.58G 6s
  7400K .......... .......... .......... .......... .......... 20% 1.74G 6s
  7450K .......... .......... .......... .......... .......... 21% 2.44G 6s
  7500K .......... .......... .......... .......... .......... 21% 2.33G 6s
  7550K .......... .......... .......... .......... .......... 21% 1.55G 6s
  7600K .......... .......... .......... .......... .......... 21% 1.00G 6s
  7650K .......... .......... .......... .......... .......... 21% 1.81G 6s
  7700K .......... .......... .......... .......... .......... 21% 2.42G 6s
  7750K .......... .......... .......... .......... .......... 21% 2.06G 6s
  7800K .......... .......... .......... .......... .......... 22% 2.01G 6s
  7850K .......... .......... .......... .......... .......... 22% 2.34G 5s
  7900K .......... .......... .......... .......... .......... 22% 1.43G 5s
  7950K .......... .......... .......... .......... .......... 22% 1.59G 5s
  8000K .......... .......... .......... .......... .......... 22% 2.50G 5s
  8050K .......... .......... .......... .......... .......... 22% 2.61G 5s
  8100K .......... .......... .......... .......... .......... 22% 2.95G 5s
  8150K .......... .......... .......... .......... .......... 23% 2.18G 5s
  8200K .......... .......... .......... .......... .......... 23% 2.59G 5s
  8250K .......... .......... .......... .......... .......... 23% 2.64G 5s
  8300K .......... .......... .......... .......... .......... 23% 2.56G 5s
  8350K .......... .......... .......... .......... .......... 23% 2.24G 5s
  8400K .......... .......... .......... .......... .......... 23% 2.71G 5s
  8450K .......... .......... .......... .......... .......... 23% 2.44G 5s
  8500K .......... .......... .......... .......... .......... 23% 2.99G 5s
  8550K .......... .......... .......... .......... .......... 24% 2.63G 5s
  8600K .......... .......... .......... .......... .......... 24% 3.18G 5s
  8650K .......... .......... .......... .......... .......... 24% 3.13G 5s
  8700K .......... .......... .......... .......... .......... 24% 3.10G 5s
  8750K .......... .......... .......... .......... .......... 24% 5.27M 5s
  8800K .......... .......... .......... .......... .......... 24%  130M 5s
  8850K .......... .......... .......... .......... .......... 24%  278M 5s
  8900K .......... .......... .......... .......... .......... 25%  460M 5s
  8950K .......... .......... .......... .......... .......... 25%  243M 5s
  9000K .......... .......... .......... .......... .......... 25%  274M 5s
  9050K .......... .......... .......... .......... .......... 25%  324M 5s
  9100K .......... .......... .......... .......... .......... 25%  571M 5s
  9150K .......... .......... .......... .......... .......... 25%  211M 5s
  9200K .......... .......... .......... .......... .......... 25%  192M 5s
  9250K .......... .......... .......... .......... .......... 26%  239M 5s
  9300K .......... .......... .......... .......... .......... 26%  557M 5s
  9350K .......... .......... .......... .......... .......... 26%  328M 5s
  9400K .......... .......... .......... .......... .......... 26%  425M 5s
  9450K .......... .......... .......... .......... .......... 26% 2.34M 5s
  9500K .......... .......... .......... .......... .......... 26% 67.3M 5s
  9550K .......... .......... .......... .......... .......... 26% 83.9M 5s
  9600K .......... .......... .......... .......... .......... 27%  509M 5s
  9650K .......... .......... .......... .......... .......... 27%  286M 5s
  9700K .......... .......... .......... .......... .......... 27%  181M 5s
  9750K .......... .......... .......... .......... .......... 27% 1.25G 5s
  9800K .......... .......... .......... .......... .......... 27% 1.76G 5s
  9850K .......... .......... .......... .......... .......... 27% 1.78G 5s
  9900K .......... .......... .......... .......... .......... 27% 1.46G 5s
  9950K .......... .......... .......... .......... .......... 28% 1.74G 5s
 10000K .......... .......... .......... .......... .......... 28% 1.97G 5s
 10050K .......... .......... .......... .......... .......... 28% 2.42G 5s
 10100K .......... .......... .......... .......... .......... 28% 2.09G 5s
 10150K .......... .......... .......... .......... .......... 28% 2.47G 5s
 10200K .......... .......... .......... .......... .......... 28% 2.50G 5s
 10250K .......... .......... .......... .......... .......... 28% 2.40G 5s
 10300K .......... .......... .......... .......... .......... 29% 2.13G 5s
 10350K .......... .......... .......... .......... .......... 29% 2.48G 4s
 10400K .......... .......... .......... .......... .......... 29% 2.47G 4s
 10450K .......... .......... .......... .......... .......... 29% 2.50G 4s
 10500K .......... .......... .......... .......... .......... 29% 1.74G 4s
 10550K .......... .......... .......... .......... .......... 29% 2.48G 4s
 10600K .......... .......... .......... .......... .......... 29% 16.6M 4s
 10650K .......... .......... .......... .......... .......... 30%  495M 4s
 10700K .......... .......... .......... .......... .......... 30%  319M 4s
 10750K .......... .......... .......... .......... .......... 30%  353M 4s
 10800K .......... .......... .......... .......... .......... 30% 1.08G 4s
 10850K .......... .......... .......... .......... .......... 30% 2.25G 4s
 10900K .......... .......... .......... .......... .......... 30%  224M 4s
 10950K .......... .......... .......... .......... .......... 30%  171M 4s
 11000K .......... .......... .......... .......... .......... 31%  729M 4s
 11050K .......... .......... .......... .......... .......... 31%  208M 4s
 11100K .......... .......... .......... .......... .......... 31% 2.69G 4s
 11150K .......... .......... .......... .......... .......... 31%  163M 4s
 11200K .......... .......... .......... .......... .......... 31%  994M 4s
 11250K .......... .......... .......... .......... .......... 31%  268M 4s
 11300K .......... .......... .......... .......... .......... 31% 2.88G 4s
 11350K .......... .......... .......... .......... .......... 31% 2.17G 4s
 11400K .......... .......... .......... .......... .......... 32% 2.29G 4s
 11450K .......... .......... .......... .......... .......... 32% 2.84G 4s
 11500K .......... .......... .......... .......... .......... 32% 12.5M 4s
 11550K .......... .......... .......... .......... .......... 32%  131M 4s
 11600K .......... .......... .......... .......... .......... 32%  200M 4s
 11650K .......... .......... .......... .......... .......... 32%  204M 4s
 11700K .......... .......... .......... .......... .......... 32%  389M 4s
 11750K .......... .......... .......... .......... .......... 33%  358M 4s
 11800K .......... .......... .......... .......... .......... 33%  586M 4s
 11850K .......... .......... .......... .......... .......... 33% 13.4M 4s
 11900K .......... .......... .......... .......... .......... 33%  248M 4s
 11950K .......... .......... .......... .......... .......... 33%  106M 4s
 12000K .......... .......... .......... .......... .......... 33%  240M 4s
 12050K .......... .......... .......... .......... .......... 33%  240M 4s
 12100K .......... .......... .......... .......... .......... 34%  284M 4s
 12150K .......... .......... .......... .......... .......... 34%  143M 4s
 12200K .......... .......... .......... .......... .......... 34%  425M 4s
 12250K .......... .......... .......... .......... .......... 34%  173M 4s
 12300K .......... .......... .......... .......... .......... 34%  318M 4s
 12350K .......... .......... .......... .......... .......... 34%  269M 4s
 12400K .......... .......... .......... .......... .......... 34%  103M 4s
 12450K .......... .......... .......... .......... .......... 35% 69.2M 4s
 12500K .......... .......... .......... .......... .......... 35% 63.5M 4s
 12550K .......... .......... .......... .......... .......... 35% 3.97M 4s
 12600K .......... .......... .......... .......... .......... 35% 76.1M 4s
 12650K .......... .......... .......... .......... .......... 35% 17.9M 4s
 12700K .......... .......... .......... .......... .......... 35%  140M 4s
 12750K .......... .......... .......... .......... .......... 35% 38.5M 4s
 12800K .......... .......... .......... .......... .......... 36% 1.77G 4s
 12850K .......... .......... .......... .......... .......... 36% 2.47G 4s
 12900K .......... .......... .......... .......... .......... 36% 2.13G 4s
 12950K .......... .......... .......... .......... .......... 36% 2.48G 4s
 13000K .......... .......... .......... .......... .......... 36% 2.50G 4s
 13050K .......... .......... .......... .......... .......... 36% 2.45G 4s
 13100K .......... .......... .......... .......... .......... 36% 1.67G 4s
 13150K .......... .......... .......... .......... .......... 37% 2.01G 4s
 13200K .......... .......... .......... .......... .......... 37% 9.63M 4s
 13250K .......... .......... .......... .......... .......... 37%  481M 4s
 13300K .......... .......... .......... .......... .......... 37%  138M 4s
 13350K .......... .......... .......... .......... .......... 37% 2.38G 4s
 13400K .......... .......... .......... .......... .......... 37%  376M 4s
 13450K .......... .......... .......... .......... .......... 37%  583M 4s
 13500K .......... .......... .......... .......... .......... 38%  136M 4s
 13550K .......... .......... .......... .......... .......... 38%  192M 4s
 13600K .......... .......... .......... .......... .......... 38%  120M 4s
 13650K .......... .......... .......... .......... .......... 38% 71.5M 4s
 13700K .......... .......... .......... .......... .......... 38%  914M 4s
 13750K .......... .......... .......... .......... .......... 38% 3.06G 3s
 13800K .......... .......... .......... .......... .......... 38% 58.2M 3s
 13850K .......... .......... .......... .......... .......... 38% 3.08G 3s
 13900K .......... .......... .......... .......... .......... 39% 3.15G 3s
 13950K .......... .......... .......... .......... .......... 39% 2.68G 3s
 14000K .......... .......... .......... .......... .......... 39% 3.15G 3s
 14050K .......... .......... .......... .......... .......... 39% 3.13G 3s
 14100K .......... .......... .......... .......... .......... 39% 3.18G 3s
 14150K .......... .......... .......... .......... .......... 39% 2.50G 3s
 14200K .......... .......... .......... .......... .......... 39% 3.15G 3s
 14250K .......... .......... .......... .......... .......... 40% 3.30G 3s
 14300K .......... .......... .......... .......... .......... 40%  143M 3s
 14350K .......... .......... .......... .......... .......... 40% 51.6M 3s
 14400K .......... .......... .......... .......... .......... 40% 41.0M 3s
 14450K .......... .......... .......... .......... .......... 40% 48.5M 3s
 14500K .......... .......... .......... .......... .......... 40% 44.3M 3s
 14550K .......... .......... .......... .......... .......... 40% 48.7M 3s
 14600K .......... .......... .......... .......... .......... 41% 47.9M 3s
 14650K .......... .......... .......... .......... .......... 41%  104M 3s
 14700K .......... .......... .......... .......... .......... 41%  188M 3s
 14750K .......... .......... .......... .......... .......... 41%  166M 3s
 14800K .......... .......... .......... .......... .......... 41%  133M 3s
 14850K .......... .......... .......... .......... .......... 41%  250M 3s
 14900K .......... .......... .......... .......... .......... 41%  162M 3s
 14950K .......... .......... .......... .......... .......... 42% 3.34M 3s
 15000K .......... .......... .......... .......... .......... 42% 92.1M 3s
 15050K .......... .......... .......... .......... .......... 42% 62.7M 3s
 15100K .......... .......... .......... .......... .......... 42% 71.3M 3s
 15150K .......... .......... .......... .......... .......... 42%  115M 3s
 15200K .......... .......... .......... .......... .......... 42% 2.08G 3s
 15250K .......... .......... .......... .......... .......... 42% 2.47G 3s
 15300K .......... .......... .......... .......... .......... 43% 2.48G 3s
 15350K .......... .......... .......... .......... .......... 43% 2.48G 3s
 15400K .......... .......... .......... .......... .......... 43% 2.16G 3s
 15450K .......... .......... .......... .......... .......... 43% 2.50G 3s
 15500K .......... .......... .......... .......... .......... 43% 2.47G 3s
 15550K .......... .......... .......... .......... .......... 43% 2.50G 3s
 15600K .......... .......... .......... .......... .......... 43% 2.16G 3s
 15650K .......... .......... .......... .......... .......... 44% 2.51G 3s
 15700K .......... .......... .......... .......... .......... 44% 6.44M 3s
 15750K .......... .......... .......... .......... .......... 44%  137M 3s
 15800K .......... .......... .......... .......... .......... 44% 2.95G 3s
 15850K .......... .......... .......... .......... .......... 44% 52.6M 3s
 15900K .......... .......... .......... .......... .......... 44% 1.94G 3s
 15950K .......... .......... .......... .......... .......... 44% 2.53G 3s
 16000K .......... .......... .......... .......... .......... 45% 2.16G 3s
 16050K .......... .......... .......... .......... .......... 45% 2.53G 3s
 16100K .......... .......... .......... .......... .......... 45% 2.47G 3s
 16150K .......... .......... .......... .......... .......... 45% 2.51G 3s
 16200K .......... .......... .......... .......... .......... 45% 2.05G 3s
 16250K .......... .......... .......... .......... .......... 45% 3.20G 3s
 16300K .......... .......... .......... .......... .......... 45% 3.18G 3s
 16350K .......... .......... .......... .......... .......... 46% 3.15G 3s
 16400K .......... .......... .......... .......... .......... 46% 2.75G 3s
 16450K .......... .......... .......... .......... .......... 46% 3.23G 3s
 16500K .......... .......... .......... .......... .......... 46% 3.44G 3s
 16550K .......... .......... .......... .......... .......... 46% 3.36G 3s
 16600K .......... .......... .......... .......... .......... 46% 37.2M 3s
 16650K .......... .......... .......... .......... .......... 46% 37.2M 3s
 16700K .......... .......... .......... .......... .......... 46% 77.0M 3s
 16750K .......... .......... .......... .......... .......... 47% 39.2M 3s
 16800K .......... .......... .......... .......... .......... 47% 50.0M 3s
 16850K .......... .......... .......... .......... .......... 47% 33.0M 3s
 16900K .......... .......... .......... .......... .......... 47% 42.6M 3s
 16950K .......... .......... .......... .......... .......... 47%  132M 3s
 17000K .......... .......... .......... .......... .......... 47%  343M 3s
 17050K .......... .......... .......... .......... .......... 47%  217M 3s
 17100K .......... .......... .......... .......... .......... 48%  185M 3s
 17150K .......... .......... .......... .......... .......... 48% 2.71M 3s
 17200K .......... .......... .......... .......... .......... 48% 1.71G 3s
 17250K .......... .......... .......... .......... .......... 48% 1.89G 3s
 17300K .......... .......... .......... .......... .......... 48% 1.74G 3s
 17350K .......... .......... .......... .......... .......... 48% 1.63G 3s
 17400K .......... .......... .......... .......... .......... 48% 1.87G 3s
 17450K .......... .......... .......... .......... .......... 49% 1.89G 3s
 17500K .......... .......... .......... .......... .......... 49% 1.85G 3s
 17550K .......... .......... .......... .......... .......... 49% 1.48G 3s
 17600K .......... .......... .......... .......... .......... 49% 2.28G 3s
 17650K .......... .......... .......... .......... .......... 49% 2.01G 3s
 17700K .......... .......... .......... .......... .......... 49% 1.73G 3s
 17750K .......... .......... .......... .......... .......... 49% 1.38G 3s
 17800K .......... .......... .......... .......... .......... 50% 1.69G 3s
 17850K .......... .......... .......... .......... .......... 50% 2.47G 3s
 17900K .......... .......... .......... .......... .......... 50% 2.63G 3s
 17950K .......... .......... .......... .......... .......... 50% 2.23G 3s
 18000K .......... .......... .......... .......... .......... 50% 18.9M 3s
 18050K .......... .......... .......... .......... .......... 50%  142M 3s
 18100K .......... .......... .......... .......... .......... 50%  265M 3s
 18150K .......... .......... .......... .......... .......... 51% 8.45M 3s
 18200K .......... .......... .......... .......... .......... 51% 69.8M 3s
 18250K .......... .......... .......... .......... .......... 51%  111M 3s
 18300K .......... .......... .......... .......... .......... 51%  331M 3s
 18350K .......... .......... .......... .......... .......... 51%  215M 3s
 18400K .......... .......... .......... .......... .......... 51% 22.7M 3s
 18450K .......... .......... .......... .......... .......... 51%  122M 3s
 18500K .......... .......... .......... .......... .......... 52%  139M 3s
 18550K .......... .......... .......... .......... .......... 52% 8.72M 3s
 18600K .......... .......... .......... .......... .......... 52% 89.4M 3s
 18650K .......... .......... .......... .......... .......... 52% 74.0M 3s
 18700K .......... .......... .......... .......... .......... 52%  134M 3s
 18750K .......... .......... .......... .......... .......... 52%  826M 3s
 18800K .......... .......... .......... .......... .......... 52% 28.2M 3s
 18850K .......... .......... .......... .......... .......... 53% 79.0M 3s
 18900K .......... .......... .......... .......... .......... 53%  125M 3s
 18950K .......... .......... .......... .......... .......... 53% 8.89M 3s
 19000K .......... .......... .......... .......... .......... 53%  119M 3s
 19050K .......... .......... .......... .......... .......... 53% 60.5M 3s
 19100K .......... .......... .......... .......... .......... 53% 62.7M 3s
 19150K .......... .......... .......... .......... .......... 53%  187M 3s
 19200K .......... .......... .......... .......... .......... 54% 71.1M 3s
 19250K .......... .......... .......... .......... .......... 54% 50.8M 3s
 19300K .......... .......... .......... .......... .......... 54%  134M 3s
 19350K .......... .......... .......... .......... .......... 54% 9.17M 3s
 19400K .......... .......... .......... .......... .......... 54% 71.9M 3s
 19450K .......... .......... .......... .......... .......... 54% 59.0M 3s
 19500K .......... .......... .......... .......... .......... 54% 52.4M 3s
 19550K .......... .......... .......... .......... .......... 54%  126M 3s
 19600K .......... .......... .......... .......... .......... 55%  128M 3s
 19650K .......... .......... .......... .......... .......... 55% 91.2M 3s
 19700K .......... .......... .......... .......... .......... 55% 58.8M 2s
 19750K .......... .......... .......... .......... .......... 55% 12.8M 3s
 19800K .......... .......... .......... .......... .......... 55% 25.7M 3s
 19850K .......... .......... .......... .......... .......... 55% 57.1M 2s
 19900K .......... .......... .......... .......... .......... 55% 39.1M 2s
 19950K .......... .......... .......... .......... .......... 56%  169M 2s
 20000K .......... .......... .......... .......... .......... 56%  160M 2s
 20050K .......... .......... .......... .......... .......... 56% 72.5M 2s
 20100K .......... .......... .......... .......... .......... 56% 73.5M 2s
 20150K .......... .......... .......... .......... .......... 56%  105M 2s
 20200K .......... .......... .......... .......... .......... 56% 9.46M 2s
 20250K .......... .......... .......... .......... .......... 56% 63.6M 2s
 20300K .......... .......... .......... .......... .......... 57% 33.9M 2s
 20350K .......... .......... .......... .......... .......... 57% 78.0M 2s
 20400K .......... .......... .......... .......... .......... 57%  129M 2s
 20450K .......... .......... .......... .......... .......... 57%  296M 2s
 20500K .......... .......... .......... .......... .......... 57% 70.2M 2s
 20550K .......... .......... .......... .......... .......... 57%  131M 2s
 20600K .......... .......... .......... .......... .......... 57% 9.30M 2s
 20650K .......... .......... .......... .......... .......... 58% 72.9M 2s
 20700K .......... .......... .......... .......... .......... 58% 89.7M 2s
 20750K .......... .......... .......... .......... .......... 58% 31.7M 2s
 20800K .......... .......... .......... .......... .......... 58% 95.5M 2s
 20850K .......... .......... .......... .......... .......... 58%  118M 2s
 20900K .......... .......... .......... .......... .......... 58%  163M 2s
 20950K .......... .......... .......... .......... .......... 58% 94.6M 2s
 21000K .......... .......... .......... .......... .......... 59% 9.59M 2s
 21050K .......... .......... .......... .......... .......... 59% 88.9M 2s
 21100K .......... .......... .......... .......... .......... 59% 60.0M 2s
 21150K .......... .......... .......... .......... .......... 59% 31.1M 2s
 21200K .......... .......... .......... .......... .......... 59%  110M 2s
 21250K .......... .......... .......... .......... .......... 59% 69.9M 2s
 21300K .......... .......... .......... .......... .......... 59%  199M 2s
 21350K .......... .......... .......... .......... .......... 60%  106M 2s
 21400K .......... .......... .......... .......... .......... 60%  144M 2s
 21450K .......... .......... .......... .......... .......... 60% 9.59M 2s
 21500K .......... .......... .......... .......... .......... 60% 44.0M 2s
 21550K .......... .......... .......... .......... .......... 60% 35.7M 2s
 21600K .......... .......... .......... .......... .......... 60% 84.4M 2s
 21650K .......... .......... .......... .......... .......... 60% 73.7M 2s
 21700K .......... .......... .......... .......... .......... 61%  132M 2s
 21750K .......... .......... .......... .......... .......... 61%  175M 2s
 21800K .......... .......... .......... .......... .......... 61%  151M 2s
 21850K .......... .......... .......... .......... .......... 61% 9.46M 2s
 21900K .......... .......... .......... .......... .......... 61% 96.6M 2s
 21950K .......... .......... .......... .......... .......... 61% 80.9M 2s
 22000K .......... .......... .......... .......... .......... 61% 32.3M 2s
 22050K .......... .......... .......... .......... .......... 62% 68.7M 2s
 22100K .......... .......... .......... .......... .......... 62% 60.9M 2s
 22150K .......... .......... .......... .......... .......... 62%  125M 2s
 22200K .......... .......... .......... .......... .......... 62%  130M 2s
 22250K .......... .......... .......... .......... .......... 62%  233M 2s
 22300K .......... .......... .......... .......... .......... 62% 9.96M 2s
 22350K .......... .......... .......... .......... .......... 62% 62.3M 2s
 22400K .......... .......... .......... .......... .......... 62% 89.5M 2s
 22450K .......... .......... .......... .......... .......... 63% 31.6M 2s
 22500K .......... .......... .......... .......... .......... 63% 58.6M 2s
 22550K .......... .......... .......... .......... .......... 63% 90.4M 2s
 22600K .......... .......... .......... .......... .......... 63%  154M 2s
 22650K .......... .......... .......... .......... .......... 63%  152M 2s
 22700K .......... .......... .......... .......... .......... 63%  152M 2s
 22750K .......... .......... .......... .......... .......... 63% 10.1M 2s
 22800K .......... .......... .......... .......... .......... 64% 46.3M 2s
 22850K .......... .......... .......... .......... .......... 64% 37.8M 2s
 22900K .......... .......... .......... .......... .......... 64% 93.4M 2s
 22950K .......... .......... .......... .......... .......... 64% 46.7M 2s
 23000K .......... .......... .......... .......... .......... 64%  134M 2s
 23050K .......... .......... .......... .......... .......... 64% 93.6M 2s
 23100K .......... .......... .......... .......... .......... 64% 83.7M 2s
 23150K .......... .......... .......... .......... .......... 65% 12.1M 2s
 23200K .......... .......... .......... .......... .......... 65% 71.9M 2s
 23250K .......... .......... .......... .......... .......... 65% 45.3M 2s
 23300K .......... .......... .......... .......... .......... 65% 36.8M 2s
 23350K .......... .......... .......... .......... .......... 65% 87.7M 2s
 23400K .......... .......... .......... .......... .......... 65% 49.3M 2s
 23450K .......... .......... .......... .......... .......... 65%  118M 2s
 23500K .......... .......... .......... .......... .......... 66%  128M 2s
 23550K .......... .......... .......... .......... .......... 66% 85.0M 2s
 23600K .......... .......... .......... .......... .......... 66% 11.9M 2s
 23650K .......... .......... .......... .......... .......... 66%  124M 2s
 23700K .......... .......... .......... .......... .......... 66% 40.7M 2s
 23750K .......... .......... .......... .......... .......... 66% 30.7M 2s
 23800K .......... .......... .......... .......... .......... 66%  150M 2s
 23850K .......... .......... .......... .......... .......... 67% 45.2M 2s
 23900K .......... .......... .......... .......... .......... 67%  166M 2s
 23950K .......... .......... .......... .......... .......... 67% 83.8M 2s
 24000K .......... .......... .......... .......... .......... 67%  122M 2s
 24050K .......... .......... .......... .......... .......... 67% 11.8M 2s
 24100K .......... .......... .......... .......... .......... 67% 80.4M 2s
 24150K .......... .......... .......... .......... .......... 67% 56.1M 2s
 24200K .......... .......... .......... .......... .......... 68% 27.6M 2s
 24250K .......... .......... .......... .......... .......... 68%  105M 2s
 24300K .......... .......... .......... .......... .......... 68% 50.6M 2s
 24350K .......... .......... .......... .......... .......... 68%  224M 2s
 24400K .......... .......... .......... .......... .......... 68% 67.5M 2s
 24450K .......... .......... .......... .......... .......... 68% 14.7M 2s
 24500K .......... .......... .......... .......... .......... 68% 46.0M 2s
 24550K .......... .......... .......... .......... .......... 69% 95.6M 2s
 24600K .......... .......... .......... .......... .......... 69% 23.4M 2s
 24650K .......... .......... .......... .......... .......... 69% 63.5M 2s
 24700K .......... .......... .......... .......... .......... 69%  204M 2s
 24750K .......... .......... .......... .......... .......... 69% 46.0M 2s
 24800K .......... .......... .......... .......... .......... 69%  136M 2s
 24850K .......... .......... .......... .......... .......... 69% 69.7M 2s
 24900K .......... .......... .......... .......... .......... 69% 14.7M 2s
 24950K .......... .......... .......... .......... .......... 70% 59.9M 2s
 25000K .......... .......... .......... .......... .......... 70%  126M 2s
 25050K .......... .......... .......... .......... .......... 70% 21.8M 2s
 25100K .......... .......... .......... .......... .......... 70% 82.0M 2s
 25150K .......... .......... .......... .......... .......... 70%  162M 2s
 25200K .......... .......... .......... .......... .......... 70% 46.0M 2s
 25250K .......... .......... .......... .......... .......... 70% 82.3M 2s
 25300K .......... .......... .......... .......... .......... 71% 76.3M 2s
 25350K .......... .......... .......... .......... .......... 71% 15.5M 2s
 25400K .......... .......... .......... .......... .......... 71% 49.3M 2s
 25450K .......... .......... .......... .......... .......... 71% 69.7M 2s
 25500K .......... .......... .......... .......... .......... 71% 26.9M 2s
 25550K .......... .......... .......... .......... .......... 71% 74.3M 2s
 25600K .......... .......... .......... .......... .......... 71% 83.1M 2s
 25650K .......... .......... .......... .......... .......... 72% 53.3M 2s
 25700K .......... .......... .......... .......... .......... 72%  100M 2s
 25750K .......... .......... .......... .......... .......... 72% 69.5M 2s
 25800K .......... .......... .......... .......... .......... 72% 15.4M 2s
 25850K .......... .......... .......... .......... .......... 72% 45.5M 2s
 25900K .......... .......... .......... .......... .......... 72% 91.9M 2s
 25950K .......... .......... .......... .......... .......... 72% 25.5M 2s
 26000K .......... .......... .......... .......... .......... 73%  156M 2s
 26050K .......... .......... .......... .......... .......... 73% 89.1M 2s
 26100K .......... .......... .......... .......... .......... 73% 39.1M 2s
 26150K .......... .......... .......... .......... .......... 73%  123M 2s
 26200K .......... .......... .......... .......... .......... 73%  115M 2s
 26250K .......... .......... .......... .......... .......... 73% 14.8M 2s
 26300K .......... .......... .......... .......... .......... 73% 49.8M 2s
 26350K .......... .......... .......... .......... .......... 74% 79.5M 2s
 26400K .......... .......... .......... .......... .......... 74% 23.6M 2s
 26450K .......... .......... .......... .......... .......... 74% 88.3M 2s
 26500K .......... .......... .......... .......... .......... 74%  111M 2s
 26550K .......... .......... .......... .......... .......... 74% 43.2M 2s
 26600K .......... .......... .......... .......... .......... 74%  106M 1s
 26650K .......... .......... .......... .......... .......... 74%  151M 1s
 26700K .......... .......... .......... .......... .......... 75% 49.9M 1s
 26750K .......... .......... .......... .......... .......... 75% 15.2M 1s
 26800K .......... .......... .......... .......... .......... 75% 69.2M 1s
 26850K .......... .......... .......... .......... .......... 75% 94.6M 1s
 26900K .......... .......... .......... .......... .......... 75% 23.7M 1s
 26950K .......... .......... .......... .......... .......... 75%  152M 1s
 27000K .......... .......... .......... .......... .......... 75% 34.9M 1s
 27050K .......... .......... .......... .......... .......... 76%  221M 1s
 27100K .......... .......... .......... .......... .......... 76% 77.7M 1s
 27150K .......... .......... .......... .......... .......... 76% 69.9M 1s
 27200K .......... .......... .......... .......... .......... 76% 15.7M 1s
 27250K .......... .......... .......... .......... .......... 76% 50.5M 1s
 27300K .......... .......... .......... .......... .......... 76% 82.0M 1s
 27350K .......... .......... .......... .......... .......... 76% 23.4M 1s
 27400K .......... .......... .......... .......... .......... 77%  172M 1s
 27450K .......... .......... .......... .......... .......... 77% 38.6M 1s
 27500K .......... .......... .......... .......... .......... 77%  104M 1s
 27550K .......... .......... .......... .......... .......... 77%  153M 1s
 27600K .......... .......... .......... .......... .......... 77% 78.4M 1s
 27650K .......... .......... .......... .......... .......... 77% 14.2M 1s
 27700K .......... .......... .......... .......... .......... 77% 64.1M 1s
 27750K .......... .......... .......... .......... .......... 77%  127M 1s
 27800K .......... .......... .......... .......... .......... 78% 19.1M 1s
 27850K .......... .......... .......... .......... .......... 78%  142M 1s
 27900K .......... .......... .......... .......... .......... 78% 38.5M 1s
 27950K .......... .......... .......... .......... .......... 78%  126M 1s
 28000K .......... .......... .......... .......... .......... 78%  323M 1s
 28050K .......... .......... .......... .......... .......... 78% 60.7M 1s
 28100K .......... .......... .......... .......... .......... 78% 14.7M 1s
 28150K .......... .......... .......... .......... .......... 79% 67.9M 1s
 28200K .......... .......... .......... .......... .......... 79% 95.3M 1s
 28250K .......... .......... .......... .......... .......... 79% 22.4M 1s
 28300K .......... .......... .......... .......... .......... 79%  132M 1s
 28350K .......... .......... .......... .......... .......... 79% 40.2M 1s
 28400K .......... .......... .......... .......... .......... 79% 72.4M 1s
 28450K .......... .......... .......... .......... .......... 79%  208M 1s
 28500K .......... .......... .......... .......... .......... 80% 80.7M 1s
 28550K .......... .......... .......... .......... .......... 80% 21.0M 1s
 28600K .......... .......... .......... .......... .......... 80% 36.8M 1s
 28650K .......... .......... .......... .......... .......... 80% 57.2M 1s
 28700K .......... .......... .......... .......... .......... 80% 21.7M 1s
 28750K .......... .......... .......... .......... .......... 80% 99.2M 1s
 28800K .......... .......... .......... .......... .......... 80% 82.3M 1s
 28850K .......... .......... .......... .......... .......... 81% 55.3M 1s
 28900K .......... .......... .......... .......... .......... 81% 77.1M 1s
 28950K .......... .......... .......... .......... .......... 81%  170M 1s
 29000K .......... .......... .......... .......... .......... 81% 20.9M 1s
 29050K .......... .......... .......... .......... .......... 81% 32.7M 1s
 29100K .......... .......... .......... .......... .......... 81% 61.3M 1s
 29150K .......... .......... .......... .......... .......... 81% 21.9M 1s
 29200K .......... .......... .......... .......... .......... 82% 78.6M 1s
 29250K .......... .......... .......... .......... .......... 82%  105M 1s
 29300K .......... .......... .......... .......... .......... 82% 67.1M 1s
 29350K .......... .......... .......... .......... .......... 82% 71.5M 1s
 29400K .......... .......... .......... .......... .......... 82%  123M 1s
 29450K .......... .......... .......... .......... .......... 82% 75.0M 1s
 29500K .......... .......... .......... .......... .......... 82% 14.5M 1s
 29550K .......... .......... .......... .......... .......... 83% 79.4M 1s
 29600K .......... .......... .......... .......... .......... 83%  100M 1s
 29650K .......... .......... .......... .......... .......... 83% 21.5M 1s
 29700K .......... .......... .......... .......... .......... 83% 75.9M 1s
 29750K .......... .......... .......... .......... .......... 83% 62.3M 1s
 29800K .......... .......... .......... .......... .......... 83% 91.6M 1s
 29850K .......... .......... .......... .......... .......... 83% 57.8M 1s
 29900K .......... .......... .......... .......... .......... 84%  123M 1s
 29950K .......... .......... .......... .......... .......... 84% 19.5M 1s
 30000K .......... .......... .......... .......... .......... 84% 40.3M 1s
 30050K .......... .......... .......... .......... .......... 84% 64.7M 1s
 30100K .......... .......... .......... .......... .......... 84% 22.4M 1s
 30150K .......... .......... .......... .......... .......... 84% 55.5M 1s
 30200K .......... .......... .......... .......... .......... 84%  231M 1s
 30250K .......... .......... .......... .......... .......... 85%  105M 1s
 30300K .......... .......... .......... .......... .......... 85% 42.6M 1s
 30350K .......... .......... .......... .......... .......... 85% 93.3M 1s
 30400K .......... .......... .......... .......... .......... 85% 93.6M 1s
 30450K .......... .......... .......... .......... .......... 85% 17.1M 1s
 30500K .......... .......... .......... .......... .......... 85% 61.4M 1s
 30550K .......... .......... .......... .......... .......... 85% 20.1M 1s
 30600K .......... .......... .......... .......... .......... 85% 71.6M 1s
 30650K .......... .......... .......... .......... .......... 86% 99.5M 1s
 30700K .......... .......... .......... .......... .......... 86%  132M 1s
 30750K .......... .......... .......... .......... .......... 86%  110M 1s
 30800K .......... .......... .......... .......... .......... 86% 41.6M 1s
 30850K .......... .......... .......... .......... .......... 86% 84.6M 1s
 30900K .......... .......... .......... .......... .......... 86% 16.7M 1s
 30950K .......... .......... .......... .......... .......... 86% 96.5M 1s
 31000K .......... .......... .......... .......... .......... 87% 52.1M 1s
 31050K .......... .......... .......... .......... .......... 87% 23.4M 1s
 31100K .......... .......... .......... .......... .......... 87% 58.1M 1s
 31150K .......... .......... .......... .......... .......... 87%  143M 1s
 31200K .......... .......... .......... .......... .......... 87%  116M 1s
 31250K .......... .......... .......... .......... .......... 87% 65.6M 1s
 31300K .......... .......... .......... .......... .......... 87% 70.6M 1s
 31350K .......... .......... .......... .......... .......... 88% 79.0M 1s
 31400K .......... .......... .......... .......... .......... 88% 16.5M 1s
 31450K .......... .......... .......... .......... .......... 88% 62.5M 1s
 31500K .......... .......... .......... .......... .......... 88% 20.8M 1s
 31550K .......... .......... .......... .......... .......... 88%  118M 1s
 31600K .......... .......... .......... .......... .......... 88% 55.5M 1s
 31650K .......... .......... .......... .......... .......... 88%  290M 1s
 31700K .......... .......... .......... .......... .......... 89% 56.5M 1s
 31750K .......... .......... .......... .......... .......... 89% 71.3M 1s
 31800K .......... .......... .......... .......... .......... 89% 68.3M 1s
 31850K .......... .......... .......... .......... .......... 89% 16.9M 1s
 31900K .......... .......... .......... .......... .......... 89%  137M 1s
 31950K .......... .......... .......... .......... .......... 89% 16.6M 1s
 32000K .......... .......... .......... .......... .......... 89%  133M 1s
 32050K .......... .......... .......... .......... .......... 90% 83.9M 1s
 32100K .......... .......... .......... .......... .......... 90% 67.1M 1s
 32150K .......... .......... .......... .......... .......... 90%  307M 1s
 32200K .......... .......... .......... .......... .......... 90% 67.9M 1s
 32250K .......... .......... .......... .......... .......... 90% 75.5M 1s
 32300K .......... .......... .......... .......... .......... 90% 15.0M 1s
 32350K .......... .......... .......... .......... .......... 90%  197M 1s
 32400K .......... .......... .......... .......... .......... 91% 69.6M 1s
 32450K .......... .......... .......... .......... .......... 91% 17.7M 1s
 32500K .......... .......... .......... .......... .......... 91%  193M 1s
 32550K .......... .......... .......... .......... .......... 91% 57.3M 1s
 32600K .......... .......... .......... .......... .......... 91%  145M 1s
 32650K .......... .......... .......... .......... .......... 91%  109M 0s
 32700K .......... .......... .......... .......... .......... 91% 55.8M 0s
 32750K .......... .......... .......... .......... .......... 92%  141M 0s
 32800K .......... .......... .......... .......... .......... 92% 14.2M 0s
 32850K .......... .......... .......... .......... .......... 92%  111M 0s
 32900K .......... .......... .......... .......... .......... 92% 16.2M 0s
 32950K .......... .......... .......... .......... .......... 92%  104M 0s
 33000K .......... .......... .......... .......... .......... 92%  279M 0s
 33050K .......... .......... .......... .......... .......... 92% 95.1M 0s
 33100K .......... .......... .......... .......... .......... 93%  171M 0s
 33150K .......... .......... .......... .......... .......... 93% 98.1M 0s
 33200K .......... .......... .......... .......... .......... 93% 70.7M 0s
 33250K .......... .......... .......... .......... .......... 93% 28.7M 0s
 33300K .......... .......... .......... .......... .......... 93% 19.2M 0s
 33350K .......... .......... .......... .......... .......... 93%  117M 0s
 33400K .......... .......... .......... .......... .......... 93% 17.5M 0s
 33450K .......... .......... .......... .......... .......... 93% 96.4M 0s
 33500K .......... .......... .......... .......... .......... 94%  178M 0s
 33550K .......... .......... .......... .......... .......... 94%  160M 0s
 33600K .......... .......... .......... .......... .......... 94% 97.2M 0s
 33650K .......... .......... .......... .......... .......... 94% 60.4M 0s
 33700K .......... .......... .......... .......... .......... 94% 98.2M 0s
 33750K .......... .......... .......... .......... .......... 94% 14.1M 0s
 33800K .......... .......... .......... .......... .......... 94% 95.2M 0s
 33850K .......... .......... .......... .......... .......... 95% 17.2M 0s
 33900K .......... .......... .......... .......... .......... 95% 87.7M 0s
 33950K .......... .......... .......... .......... .......... 95% 43.4M 0s
 34000K .......... .......... .......... .......... .......... 95%  627M 0s
 34050K .......... .......... .......... .......... .......... 95%  282M 0s
 34100K .......... .......... .......... .......... .......... 95%  313M 0s
 34150K .......... .......... .......... .......... .......... 95% 66.6M 0s
 34200K .......... .......... .......... .......... .......... 96% 30.2M 0s
 34250K .......... .......... .......... .......... .......... 96% 20.1M 0s
 34300K .......... .......... .......... .......... .......... 96% 86.4M 0s
 34350K .......... .......... .......... .......... .......... 96% 18.2M 0s
 34400K .......... .......... .......... .......... .......... 96% 68.7M 0s
 34450K .......... .......... .......... .......... .......... 96% 47.1M 0s
 34500K .......... .......... .......... .......... .......... 96%  161M 0s
 34550K .......... .......... .......... .......... .......... 97%  385M 0s
 34600K .......... .......... .......... .......... .......... 97%  198M 0s
 34650K .......... .......... .......... .......... .......... 97%  195M 0s
 34700K .......... .......... .......... .......... .......... 97% 12.9M 0s
 34750K .......... .......... .......... .......... .......... 97%  121M 0s
 34800K .......... .......... .......... .......... .......... 97% 16.8M 0s
 34850K .......... .......... .......... .......... .......... 97%  126M 0s
 34900K .......... .......... .......... .......... .......... 98% 36.3M 0s
 34950K .......... .......... .......... .......... .......... 98% 87.5M 0s
 35000K .......... .......... .......... .......... .......... 98%  106M 0s
 35050K .......... .......... .......... .......... .......... 98%  504M 0s
 35100K .......... .......... .......... .......... .......... 98%  165M 0s
 35150K .......... .......... .......... .......... .......... 98%  143M 0s
 35200K .......... .......... .......... .......... .......... 98% 14.5M 0s
 35250K .......... .......... .......... .......... .......... 99%  143M 0s
 35300K .......... .......... .......... .......... .......... 99% 17.1M 0s
 35350K .......... .......... .......... .......... .......... 99%  102M 0s
 35400K .......... .......... .......... .......... .......... 99% 30.6M 0s
 35450K .......... .......... .......... .......... .......... 99%  101M 0s
 35500K .......... .......... .......... .......... .......... 99%  315M 0s
 35550K .......... .......... .......... .......... .......... 99% 85.6M 0s
 35600K .......... .......... .......... .......... ...       100% 1.16G=6.0s

2020-03-02 03:23:53 (48.4 Mb/s) - ‘/dev/null’ saved [36499294/36499294]

