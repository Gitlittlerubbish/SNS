--2020-02-25 22:12:37--  http://www.marn.gob.sv/inema2017.pdf%0D
Resolving www.marn.gob.sv (www.marn.gob.sv)... 104.210.5.96
Connecting to www.marn.gob.sv (www.marn.gob.sv)|104.210.5.96|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:12:37 ERROR 404: Not Found.

--2020-02-25 22:13:21--  http://www.marn.gob.sv/inema2017.pdf%0D
Resolving www.marn.gob.sv (www.marn.gob.sv)... 104.210.5.96
Connecting to www.marn.gob.sv (www.marn.gob.sv)|104.210.5.96|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:21 ERROR 404: Not Found.

