--2020-02-25 22:12:31--  http://www.transparenciafiscal.gob.sv/downloads/pdf/DC5544_CAP_21.pdf%0D
Resolving www.transparenciafiscal.gob.sv (www.transparenciafiscal.gob.sv)... 190.5.131.23, 190.57.24.31
Connecting to www.transparenciafiscal.gob.sv (www.transparenciafiscal.gob.sv)|190.5.131.23|:80... connected.
HTTP request sent, awaiting response... 302 Found
Location: http://www.transparenciafiscal.gob.sv/ptf/es/index.html [following]
--2020-02-25 22:12:31--  http://www.transparenciafiscal.gob.sv/ptf/es/index.html
Reusing existing connection to www.transparenciafiscal.gob.sv:80.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K ....                                                   18.0M=0.002s

2020-02-25 22:12:32 (18.0 Mb/s) - ‘/dev/null’ saved [4388]

--2020-02-25 22:12:32--  http://www.transparenciafiscal.gob.sv/downloads/pdf/DC5544_CAP_21.pdf%0D
Resolving www.transparenciafiscal.gob.sv (www.transparenciafiscal.gob.sv)... 190.5.131.23, 190.57.24.31
Connecting to www.transparenciafiscal.gob.sv (www.transparenciafiscal.gob.sv)|190.5.131.23|:80... connected.
HTTP request sent, awaiting response... 302 Found
Location: http://www.transparenciafiscal.gob.sv/ptf/es/index.html [following]
--2020-02-25 22:12:32--  http://www.transparenciafiscal.gob.sv/ptf/es/index.html
Reusing existing connection to www.transparenciafiscal.gob.sv:80.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K ....                                                   17.9M=0.002s

2020-02-25 22:12:32 (17.9 Mb/s) - ‘/dev/null’ saved [4388]

--2020-02-25 22:13:15--  http://www.transparenciafiscal.gob.sv/downloads/pdf/DC5544_CAP_21.pdf%0D
Resolving www.transparenciafiscal.gob.sv (www.transparenciafiscal.gob.sv)... 190.57.24.31, 190.5.131.23
Connecting to www.transparenciafiscal.gob.sv (www.transparenciafiscal.gob.sv)|190.57.24.31|:80... connected.
HTTP request sent, awaiting response... 302 Found
Location: http://www.transparenciafiscal.gob.sv/ptf/es/index.html [following]
--2020-02-25 22:13:15--  http://www.transparenciafiscal.gob.sv/ptf/es/index.html
Reusing existing connection to www.transparenciafiscal.gob.sv:80.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K ....                                                   22.5M=0.002s

2020-02-25 22:13:16 (22.5 Mb/s) - ‘/dev/null’ saved [4388]

--2020-02-25 22:13:16--  http://www.transparenciafiscal.gob.sv/downloads/pdf/DC5544_CAP_21.pdf%0D
Resolving www.transparenciafiscal.gob.sv (www.transparenciafiscal.gob.sv)... 190.57.24.31, 190.5.131.23
Connecting to www.transparenciafiscal.gob.sv (www.transparenciafiscal.gob.sv)|190.57.24.31|:80... connected.
HTTP request sent, awaiting response... 302 Found
Location: http://www.transparenciafiscal.gob.sv/ptf/es/index.html [following]
--2020-02-25 22:13:16--  http://www.transparenciafiscal.gob.sv/ptf/es/index.html
Reusing existing connection to www.transparenciafiscal.gob.sv:80.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K ....                                                   20.3M=0.002s

2020-02-25 22:13:16 (20.3 Mb/s) - ‘/dev/null’ saved [4388]

