--2020-03-02 03:25:12--  http://www.grupoacc.com.sv/Files/DEC_160.pdf
Resolving www.grupoacc.com.sv (www.grupoacc.com.sv)... 192.185.148.210
Connecting to www.grupoacc.com.sv (www.grupoacc.com.sv)|192.185.148.210|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 1707510 (1.6M) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  2% 1.66M 8s
    50K .......... .......... .......... .......... ..........  5% 3.34M 6s
   100K .......... .......... .......... .......... ..........  8%  129M 4s
   150K .......... .......... .......... .......... .......... 11% 29.3M 3s
   200K .......... .......... .......... .......... .......... 14% 3.75M 3s
   250K .......... .......... .......... .......... .......... 17% 32.4M 2s
   300K .......... .......... .......... .......... .......... 20% 3.74M 2s
   350K .......... .......... .......... .......... .......... 23%  212M 2s
   400K .......... .......... .......... .......... .......... 26% 80.3M 2s
   450K .......... .......... .......... .......... .......... 29%  180M 1s
   500K .......... .......... .......... .......... .......... 32% 59.4M 1s
   550K .......... .......... .......... .......... .......... 35% 3.70M 1s
   600K .......... .......... .......... .......... .......... 38%  309M 1s
   650K .......... .......... .......... .......... .......... 41%  109M 1s
   700K .......... .......... .......... .......... .......... 44%  104M 1s
   750K .......... .......... .......... .......... .......... 47% 84.8M 1s
   800K .......... .......... .......... .......... .......... 50% 3.67M 1s
   850K .......... .......... .......... .......... .......... 53%  203M 1s
   900K .......... .......... .......... .......... .......... 56%  463M 1s
   950K .......... .......... .......... .......... .......... 59%  243M 1s
  1000K .......... .......... .......... .......... .......... 62%  452M 1s
  1050K .......... .......... .......... .......... .......... 65%  217M 0s
  1100K .......... .......... .......... .......... .......... 68%  303M 0s
  1150K .......... .......... .......... .......... .......... 71%  144M 0s
  1200K .......... .......... .......... .......... .......... 74% 3.98M 0s
  1250K .......... .......... .......... .......... .......... 77% 45.3M 0s
  1300K .......... .......... .......... .......... .......... 80%  127M 0s
  1350K .......... .......... .......... .......... .......... 83%  128M 0s
  1400K .......... .......... .......... .......... .......... 86%  102M 0s
  1450K .......... .......... .......... .......... .......... 89%  249M 0s
  1500K .......... .......... .......... .......... .......... 92%  519M 0s
  1550K .......... .......... .......... .......... .......... 95%  374M 0s
  1600K .......... .......... .......... .......... .......... 98%  235M 0s
  1650K .......... .......                                    100%  412M=1.0s

2020-03-02 03:25:15 (13.5 Mb/s) - ‘/dev/null’ saved [1707510/1707510]

