--2020-02-25 22:14:14--  http://tecnobodega.com.sv/images/Productos/20170620311528_V7S36LA.pdf%0D
Resolving tecnobodega.com.sv (tecnobodega.com.sv)... 168.243.50.98
Connecting to tecnobodega.com.sv (tecnobodega.com.sv)|168.243.50.98|:80... connected.
HTTP request sent, awaiting response... 400 Bad Request
2020-02-25 22:14:14 ERROR 400: Bad Request.

--2020-02-25 22:14:38--  http://tecnobodega.com.sv/images/Productos/20170620311528_V7S36LA.pdf%0D
Resolving tecnobodega.com.sv (tecnobodega.com.sv)... 168.243.50.98
Connecting to tecnobodega.com.sv (tecnobodega.com.sv)|168.243.50.98|:80... connected.
HTTP request sent, awaiting response... 400 Bad Request
2020-02-25 22:14:39 ERROR 400: Bad Request.

