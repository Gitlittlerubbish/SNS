--2020-02-25 22:14:21--  https://www.diariooficial.gob.sv/diarios/do-2017/04-abril/26-04-2017.pdf%0D
Resolving www.diariooficial.gob.sv (www.diariooficial.gob.sv)... 190.86.209.40
Connecting to www.diariooficial.gob.sv (www.diariooficial.gob.sv)|190.86.209.40|:443... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:21 ERROR 404: Not Found.

--2020-02-25 22:14:40--  https://www.diariooficial.gob.sv/diarios/do-2017/04-abril/26-04-2017.pdf%0D
Resolving www.diariooficial.gob.sv (www.diariooficial.gob.sv)... 190.86.209.40
Connecting to www.diariooficial.gob.sv (www.diariooficial.gob.sv)|190.86.209.40|:443... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:41 ERROR 404: Not Found.

