--2020-02-25 22:13:45--  https://ovisss.isss.gob.sv/documentos_ofivi/Calendario_OVISSS_2020.pdf%0D
Resolving ovisss.isss.gob.sv (ovisss.isss.gob.sv)... 129.158.125.97
Connecting to ovisss.isss.gob.sv (ovisss.isss.gob.sv)|129.158.125.97|:443... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:45 ERROR 404: Not Found.

--2020-02-25 22:14:15--  https://ovisss.isss.gob.sv/documentos_ofivi/Calendario_OVISSS_2020.pdf%0D
Resolving ovisss.isss.gob.sv (ovisss.isss.gob.sv)... 129.158.125.97
Connecting to ovisss.isss.gob.sv (ovisss.isss.gob.sv)|129.158.125.97|:443... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:16 ERROR 404: Not Found.

