--2020-03-02 03:24:18--  http://www.fomilenioii.gob.sv/asset/documents/90
Resolving www.fomilenioii.gob.sv (www.fomilenioii.gob.sv)... 138.201.55.180
Connecting to www.fomilenioii.gob.sv (www.fomilenioii.gob.sv)|138.201.55.180|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: https://www.fomilenioii.gob.sv/asset/documents/90 [following]
--2020-03-02 03:24:18--  https://www.fomilenioii.gob.sv/asset/documents/90
Connecting to www.fomilenioii.gob.sv (www.fomilenioii.gob.sv)|138.201.55.180|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [application/x-download]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 7.78M
    50K .......... .......... .......... .......... .......... 17.7M
   100K .......... .......... .......... .......... ..........  124M
   150K .......... .......... .......... .......... .......... 27.0M
   200K .......... .......... .......... .......... .......... 52.0M
   250K .......... .......... .......... .......... .......... 81.1M
   300K .......... .......... .......... .......... .......... 29.8M
   350K .......... .......... .......... .......... ..........  102M
   400K .......... .......... .......... .......... .......... 91.4M
   450K .......... .......... .                                72.1M=0.1s

2020-03-02 03:24:18 (29.3 Mb/s) - ‘/dev/null’ saved [482980]

