--2020-02-25 22:12:35--  http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D419%0D
Resolving biblioteca.inu.edu.sv (biblioteca.inu.edu.sv)... 78.47.62.221
Connecting to biblioteca.inu.edu.sv (biblioteca.inu.edu.sv)|78.47.62.221|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D419/ [following]
--2020-02-25 22:12:35--  http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D419/
Reusing existing connection to biblioteca.inu.edu.sv:80.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 2.99M
    50K .......... .......... .......... .......... .......... 3.15M
   100K .......... ....                                        25.3M=0.3s

2020-02-25 22:12:36 (3.46 Mb/s) - ‘/dev/null’ saved [117408]

--2020-02-25 22:12:36--  http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D419%0D
Resolving biblioteca.inu.edu.sv (biblioteca.inu.edu.sv)... 78.47.62.221
Connecting to biblioteca.inu.edu.sv (biblioteca.inu.edu.sv)|78.47.62.221|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D419/ [following]
--2020-02-25 22:12:36--  http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D419/
Reusing existing connection to biblioteca.inu.edu.sv:80.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 2.93M
    50K .......... .......... .......... .......... .......... 4.71M
   100K .......... ....                                        14.4M=0.2s

2020-02-25 22:12:36 (3.99 Mb/s) - ‘/dev/null’ saved [117408]

--2020-02-25 22:12:36--  http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D387%0D
Resolving biblioteca.inu.edu.sv (biblioteca.inu.edu.sv)... 78.47.62.221
Connecting to biblioteca.inu.edu.sv (biblioteca.inu.edu.sv)|78.47.62.221|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D387/ [following]
--2020-02-25 22:12:36--  http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D387/
Reusing existing connection to biblioteca.inu.edu.sv:80.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 4.35M
    50K .......... .......... .......... .......... .......... 4.28M
   100K .......... ....                                        39.5M=0.2s

2020-02-25 22:12:37 (4.87 Mb/s) - ‘/dev/null’ saved [117408]

--2020-02-25 22:12:37--  http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D387%0D
Resolving biblioteca.inu.edu.sv (biblioteca.inu.edu.sv)... 78.47.62.221
Connecting to biblioteca.inu.edu.sv (biblioteca.inu.edu.sv)|78.47.62.221|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D387/ [following]
--2020-02-25 22:12:37--  http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D387/
Reusing existing connection to biblioteca.inu.edu.sv:80.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 3.36M
    50K .......... .......... .......... .......... .......... 3.83M
   100K .......... ....                                        27.8M=0.2s

2020-02-25 22:12:37 (4.03 Mb/s) - ‘/dev/null’ saved [117408]

--2020-02-25 22:13:19--  http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D419%0D
Resolving biblioteca.inu.edu.sv (biblioteca.inu.edu.sv)... 78.47.62.221
Connecting to biblioteca.inu.edu.sv (biblioteca.inu.edu.sv)|78.47.62.221|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D419/ [following]
--2020-02-25 22:13:19--  http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D419/
Reusing existing connection to biblioteca.inu.edu.sv:80.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 2.88M
    50K .......... .......... .......... .......... .......... 4.77M
   100K .......... ....                                        19.0M=0.2s

2020-02-25 22:13:19 (4.00 Mb/s) - ‘/dev/null’ saved [117408]

--2020-02-25 22:13:19--  http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D419%0D
Resolving biblioteca.inu.edu.sv (biblioteca.inu.edu.sv)... 78.47.62.221
Connecting to biblioteca.inu.edu.sv (biblioteca.inu.edu.sv)|78.47.62.221|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D419/ [following]
--2020-02-25 22:13:19--  http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D419/
Reusing existing connection to biblioteca.inu.edu.sv:80.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 4.28M
    50K .......... .......... .......... .......... .......... 3.42M
   100K .......... ....                                        26.6M=0.2s

2020-02-25 22:13:20 (4.27 Mb/s) - ‘/dev/null’ saved [117408]

--2020-02-25 22:13:20--  http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D387%0D
Resolving biblioteca.inu.edu.sv (biblioteca.inu.edu.sv)... 78.47.62.221
Connecting to biblioteca.inu.edu.sv (biblioteca.inu.edu.sv)|78.47.62.221|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D387/ [following]
--2020-02-25 22:13:20--  http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D387/
Reusing existing connection to biblioteca.inu.edu.sv:80.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 2.68M
    50K .......... .......... .......... .......... .......... 4.01M
   100K .......... ....                                        26.6M=0.3s

2020-02-25 22:13:20 (3.62 Mb/s) - ‘/dev/null’ saved [117408]

--2020-02-25 22:13:20--  http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D387%0D
Resolving biblioteca.inu.edu.sv (biblioteca.inu.edu.sv)... 78.47.62.221
Connecting to biblioteca.inu.edu.sv (biblioteca.inu.edu.sv)|78.47.62.221|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D387/ [following]
--2020-02-25 22:13:20--  http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D387/
Reusing existing connection to biblioteca.inu.edu.sv:80.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 3.41M
    50K .......... .......... .......... .......... .......... 3.45M
   100K .......... ....                                        26.2M=0.2s

2020-02-25 22:13:21 (3.86 Mb/s) - ‘/dev/null’ saved [117408]

