--2020-02-25 22:13:45--  https://www.salud.gob.sv/archivos/vigi_epide2019/Calendario_Epidemiologico_2019.pdf%0D
Resolving www.salud.gob.sv (www.salud.gob.sv)... 190.86.223.123
Connecting to www.salud.gob.sv (www.salud.gob.sv)|190.86.223.123|:443... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:48 ERROR 404: Not Found.

--2020-02-25 22:14:16--  https://www.salud.gob.sv/archivos/vigi_epide2019/Calendario_Epidemiologico_2019.pdf%0D
Resolving www.salud.gob.sv (www.salud.gob.sv)... 190.86.223.123
Connecting to www.salud.gob.sv (www.salud.gob.sv)|190.86.223.123|:443... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:18 ERROR 404: Not Found.

