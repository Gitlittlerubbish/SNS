--2020-02-25 22:12:47--  http://www.alges.org.sv/asset/documents/555%0D
Resolving www.alges.org.sv (www.alges.org.sv)... 46.4.127.171
Connecting to www.alges.org.sv (www.alges.org.sv)|46.4.127.171|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... ..........                       10.2M=0.02s

2020-02-25 22:12:48 (10.2 Mb/s) - ‘/dev/null’ saved [30726]

--2020-02-25 22:12:48--  http://www.alges.org.sv/asset/documents/555%0D
Resolving www.alges.org.sv (www.alges.org.sv)... 46.4.127.171
Connecting to www.alges.org.sv (www.alges.org.sv)|46.4.127.171|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... ..........                       10.1M=0.02s

2020-02-25 22:12:48 (10.1 Mb/s) - ‘/dev/null’ saved [30726]

--2020-02-25 22:13:25--  http://www.alges.org.sv/asset/documents/555%0D
Resolving www.alges.org.sv (www.alges.org.sv)... 46.4.127.171
Connecting to www.alges.org.sv (www.alges.org.sv)|46.4.127.171|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... ..........                       10.0M=0.02s

2020-02-25 22:13:25 (10.0 Mb/s) - ‘/dev/null’ saved [30726]

--2020-02-25 22:13:25--  http://www.alges.org.sv/asset/documents/555%0D
Resolving www.alges.org.sv (www.alges.org.sv)... 46.4.127.171
Connecting to www.alges.org.sv (www.alges.org.sv)|46.4.127.171|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... ..........                       10.0M=0.02s

2020-02-25 22:13:25 (10.0 Mb/s) - ‘/dev/null’ saved [30726]

