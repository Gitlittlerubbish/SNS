--2020-02-25 22:13:49--  https://www.isdemu.gob.sv/phocadownload/RVLV_documentos2016/ISDEMU_Guia_lectura_LEIV_con_enfoque_psicosocial.pdf%0D
Resolving www.isdemu.gob.sv (www.isdemu.gob.sv)... 72.46.153.202
Connecting to www.isdemu.gob.sv (www.isdemu.gob.sv)|72.46.153.202|:443... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:50 ERROR 404: Not Found.

--2020-02-25 22:14:19--  https://www.isdemu.gob.sv/phocadownload/RVLV_documentos2016/ISDEMU_Guia_lectura_LEIV_con_enfoque_psicosocial.pdf%0D
Resolving www.isdemu.gob.sv (www.isdemu.gob.sv)... 72.46.153.202
Connecting to www.isdemu.gob.sv (www.isdemu.gob.sv)|72.46.153.202|:443... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:19 ERROR 404: Not Found.

