--2020-02-25 22:12:59--  http://www.ute.gob.sv/publicaciones/0002.pdf%0D
Resolving www.ute.gob.sv (www.ute.gob.sv)... 190.86.186.18
Connecting to www.ute.gob.sv (www.ute.gob.sv)|190.86.186.18|:80... connected.
HTTP request sent, awaiting response... 403 Forbidden
2020-02-25 22:12:59 ERROR 403: Forbidden.

--2020-02-25 22:13:34--  http://www.ute.gob.sv/publicaciones/0002.pdf%0D
Resolving www.ute.gob.sv (www.ute.gob.sv)... 190.86.186.18
Connecting to www.ute.gob.sv (www.ute.gob.sv)|190.86.186.18|:80... connected.
HTTP request sent, awaiting response... 403 Forbidden
2020-02-25 22:13:34 ERROR 403: Forbidden.

