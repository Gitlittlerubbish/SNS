--2020-03-02 03:26:08--  http://www.isdemu.gob.sv/phocadownload/RVLV_documentos2016/ISDEMU_Guia_lectura_LEIV_con_enfoque_psicosocial.pdf
Resolving www.isdemu.gob.sv (www.isdemu.gob.sv)... 72.46.153.202
Connecting to www.isdemu.gob.sv (www.isdemu.gob.sv)|72.46.153.202|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 7185919 (6.9M) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  0% 1.45M 39s
    50K .......... .......... .......... .......... ..........  1% 2.91M 29s
   100K .......... .......... .......... .......... ..........  2% 2.87M 26s
   150K .......... .......... .......... .......... ..........  2% 3.02M 24s
   200K .......... .......... .......... .......... ..........  3% 68.4M 19s
   250K .......... .......... .......... .......... ..........  4% 3.05M 19s
   300K .......... .......... .......... .......... ..........  4% 58.1M 16s
   350K .......... .......... .......... .......... ..........  5% 3.17M 16s
   400K .......... .......... .......... .......... ..........  6%  105M 14s
   450K .......... .......... .......... .......... ..........  7%  189M 13s
   500K .......... .......... .......... .......... ..........  7% 63.3M 12s
   550K .......... .......... .......... .......... ..........  8% 3.19M 12s
   600K .......... .......... .......... .......... ..........  9%  117M 11s
   650K .......... .......... .......... .......... ..........  9%  103M 10s
   700K .......... .......... .......... .......... .......... 10% 87.7M 9s
   750K .......... .......... .......... .......... .......... 11% 53.2M 9s
   800K .......... .......... .......... .......... .......... 12% 3.40M 9s
   850K .......... .......... .......... .......... .......... 12%  126M 9s
   900K .......... .......... .......... .......... .......... 13%  140M 8s
   950K .......... .......... .......... .......... .......... 14%  134M 8s
  1000K .......... .......... .......... .......... .......... 14% 69.2M 7s
  1050K .......... .......... .......... .......... .......... 15%  214M 7s
  1100K .......... .......... .......... .......... .......... 16%  136M 7s
  1150K .......... .......... .......... .......... .......... 17% 4.00M 7s
  1200K .......... .......... .......... .......... .......... 17% 20.5M 6s
  1250K .......... .......... .......... .......... .......... 18% 86.2M 6s
  1300K .......... .......... .......... .......... .......... 19%  129M 6s
  1350K .......... .......... .......... .......... .......... 19%  106M 6s
  1400K .......... .......... .......... .......... .......... 20%  139M 5s
  1450K .......... .......... .......... .......... .......... 21% 23.2M 5s
  1500K .......... .......... .......... .......... .......... 22% 85.1M 5s
  1550K .......... .......... .......... .......... .......... 22%  382M 5s
  1600K .......... .......... .......... .......... .......... 23%  477M 5s
  1650K .......... .......... .......... .......... .......... 24% 4.23M 5s
  1700K .......... .......... .......... .......... .......... 24%  154M 5s
  1750K .......... .......... .......... .......... .......... 25%  131M 4s
  1800K .......... .......... .......... .......... .......... 26% 66.1M 4s
  1850K .......... .......... .......... .......... .......... 27%  150M 4s
  1900K .......... .......... .......... .......... .......... 27%  182M 4s
  1950K .......... .......... .......... .......... .......... 28% 83.6M 4s
  2000K .......... .......... .......... .......... .......... 29%  114M 4s
  2050K .......... .......... .......... .......... .......... 29%  100M 4s
  2100K .......... .......... .......... .......... .......... 30%  135M 4s
  2150K .......... .......... .......... .......... .......... 31% 61.5M 3s
  2200K .......... .......... .......... .......... .......... 32% 91.7M 3s
  2250K .......... .......... .......... .......... .......... 32%  136M 3s
  2300K .......... .......... .......... .......... .......... 33%  204M 3s
  2350K .......... .......... .......... .......... .......... 34% 4.41M 3s
  2400K .......... .......... .......... .......... .......... 34% 65.8M 3s
  2450K .......... .......... .......... .......... .......... 35%  354M 3s
  2500K .......... .......... .......... .......... .......... 36%  186M 3s
  2550K .......... .......... .......... .......... .......... 37%  257M 3s
  2600K .......... .......... .......... .......... .......... 37%  115M 3s
  2650K .......... .......... .......... .......... .......... 38%  126M 3s
  2700K .......... .......... .......... .......... .......... 39% 95.9M 3s
  2750K .......... .......... .......... .......... .......... 39%  200M 3s
  2800K .......... .......... .......... .......... .......... 40% 45.4M 3s
  2850K .......... .......... .......... .......... .......... 41%  204M 2s
  2900K .......... .......... .......... .......... .......... 42%  217M 2s
  2950K .......... .......... .......... .......... .......... 42%  132M 2s
  3000K .......... .......... .......... .......... .......... 43%  102M 2s
  3050K .......... .......... .......... .......... .......... 44%  101M 2s
  3100K .......... .......... .......... .......... .......... 44%  348M 2s
  3150K .......... .......... .......... .......... .......... 45% 4.47M 2s
  3200K .......... .......... .......... .......... .......... 46% 83.1M 2s
  3250K .......... .......... .......... .......... .......... 47% 95.6M 2s
  3300K .......... .......... .......... .......... .......... 47%  198M 2s
  3350K .......... .......... .......... .......... .......... 48%  188M 2s
  3400K .......... .......... .......... .......... .......... 49%  160M 2s
  3450K .......... .......... .......... .......... .......... 49%  321M 2s
  3500K .......... .......... .......... .......... .......... 50%  234M 2s
  3550K .......... .......... .......... .......... .......... 51% 97.2M 2s
  3600K .......... .......... .......... .......... .......... 52%  213M 2s
  3650K .......... .......... .......... .......... .......... 52% 46.2M 2s
  3700K .......... .......... .......... .......... .......... 53% 92.6M 2s
  3750K .......... .......... .......... .......... .......... 54%  513M 2s
  3800K .......... .......... .......... .......... .......... 54%  483M 2s
  3850K .......... .......... .......... .......... .......... 55%  193M 1s
  3900K .......... .......... .......... .......... .......... 56%  236M 1s
  3950K .......... .......... .......... .......... .......... 57% 70.0M 1s
  4000K .......... .......... .......... .......... .......... 57%  266M 1s
  4050K .......... .......... .......... .......... .......... 58% 4.67M 1s
  4100K .......... .......... .......... .......... .......... 59% 56.3M 1s
  4150K .......... .......... .......... .......... .......... 59%  131M 1s
  4200K .......... .......... .......... .......... .......... 60%  118M 1s
  4250K .......... .......... .......... .......... .......... 61%  151M 1s
  4300K .......... .......... .......... .......... .......... 61%  132M 1s
  4350K .......... .......... .......... .......... .......... 62%  117M 1s
  4400K .......... .......... .......... .......... .......... 63%  402M 1s
  4450K .......... .......... .......... .......... .......... 64%  140M 1s
  4500K .......... .......... .......... .......... .......... 64%  139M 1s
  4550K .......... .......... .......... .......... .......... 65%  309M 1s
  4600K .......... .......... .......... .......... .......... 66%  103M 1s
  4650K .......... .......... .......... .......... .......... 66%  180M 1s
  4700K .......... .......... .......... .......... .......... 67% 84.2M 1s
  4750K .......... .......... .......... .......... .......... 68%  251M 1s
  4800K .......... .......... .......... .......... .......... 69%  139M 1s
  4850K .......... .......... .......... .......... .......... 69%  390M 1s
  4900K .......... .......... .......... .......... .......... 70%  140M 1s
  4950K .......... .......... .......... .......... .......... 71% 33.4M 1s
  5000K .......... .......... .......... .......... .......... 71%  257M 1s
  5050K .......... .......... .......... .......... .......... 72% 5.99M 1s
  5100K .......... .......... .......... .......... .......... 73% 41.1M 1s
  5150K .......... .......... .......... .......... .......... 74% 60.8M 1s
  5200K .......... .......... .......... .......... .......... 74%  177M 1s
  5250K .......... .......... .......... .......... .......... 75%  103M 1s
  5300K .......... .......... .......... .......... .......... 76%  278M 1s
  5350K .......... .......... .......... .......... .......... 76%  180M 1s
  5400K .......... .......... .......... .......... .......... 77%  126M 1s
  5450K .......... .......... .......... .......... .......... 78%  235M 1s
  5500K .......... .......... .......... .......... .......... 79% 80.4M 1s
  5550K .......... .......... .......... .......... .......... 79%  134M 1s
  5600K .......... .......... .......... .......... .......... 80%  438M 1s
  5650K .......... .......... .......... .......... .......... 81%  196M 0s
  5700K .......... .......... .......... .......... .......... 81%  166M 0s
  5750K .......... .......... .......... .......... .......... 82%  166M 0s
  5800K .......... .......... .......... .......... .......... 83%  190M 0s
  5850K .......... .......... .......... .......... .......... 84%  140M 0s
  5900K .......... .......... .......... .......... .......... 84%  140M 0s
  5950K .......... .......... .......... .......... .......... 85%  201M 0s
  6000K .......... .......... .......... .......... .......... 86%  349M 0s
  6050K .......... .......... .......... .......... .......... 86%  303M 0s
  6100K .......... .......... .......... .......... .......... 87% 32.6M 0s
  6150K .......... .......... .......... .......... .......... 88% 7.05M 0s
  6200K .......... .......... .......... .......... .......... 89% 26.7M 0s
  6250K .......... .......... .......... .......... .......... 89%  123M 0s
  6300K .......... .......... .......... .......... .......... 90% 43.7M 0s
  6350K .......... .......... .......... .......... .......... 91%  108M 0s
  6400K .......... .......... .......... .......... .......... 91% 2.48G 0s
  6450K .......... .......... .......... .......... .......... 92%  118M 0s
  6500K .......... .......... .......... .......... .......... 93%  288M 0s
  6550K .......... .......... .......... .......... .......... 94%  220M 0s
  6600K .......... .......... .......... .......... .......... 94%  136M 0s
  6650K .......... .......... .......... .......... .......... 95%  516M 0s
  6700K .......... .......... .......... .......... .......... 96% 97.5M 0s
  6750K .......... .......... .......... .......... .......... 96%  161M 0s
  6800K .......... .......... .......... .......... .......... 97% 75.9M 0s
  6850K .......... .......... .......... .......... .......... 98%  408M 0s
  6900K .......... .......... .......... .......... .......... 99%  312M 0s
  6950K .......... .......... .......... .......... .......... 99%  188M 0s
  7000K .......... .......                                    100% 97.8M=2.3s

2020-03-02 03:26:11 (25.2 Mb/s) - ‘/dev/null’ saved [7185919/7185919]

