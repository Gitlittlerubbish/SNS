--2020-03-02 03:27:27--  http://www.csj.gob.sv/INV_PROF/INV_PROF/TRAMITE_AA_22_11_12.pdf
Resolving www.csj.gob.sv (www.csj.gob.sv)... 200.31.169.70
Connecting to www.csj.gob.sv (www.csj.gob.sv)|200.31.169.70|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 951003 (929K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  5% 1.02M 7s
    50K .......... .......... .......... .......... .......... 10% 2.95M 4s
   100K .......... .......... .......... .......... .......... 16%  267M 3s
   150K .......... .......... .......... .......... .......... 21% 3.06M 2s
   200K .......... .......... .......... .......... .......... 26%  217M 2s
   250K .......... .......... .......... .......... .......... 32% 3.06M 2s
   300K .......... .......... .......... .......... .......... 37%  133M 1s
   350K .......... .......... .......... .......... .......... 43%  515M 1s
   400K .......... .......... .......... .......... .......... 48% 3.21M 1s
   450K .......... .......... .......... .......... .......... 53%  116M 1s
   500K .......... .......... .......... .......... .......... 59% 80.9M 1s
   550K .......... .......... .......... .......... .......... 64%  457M 1s
   600K .......... .......... .......... .......... .......... 69%  198M 0s
   650K .......... .......... .......... .......... .......... 75% 3.39M 0s
   700K .......... .......... .......... .......... .......... 80% 98.1M 0s
   750K .......... .......... .......... .......... .......... 86%  265M 0s
   800K .......... .......... .......... .......... .......... 91% 77.9M 0s
   850K .......... .......... .......... .......... .......... 96%  152M 0s
   900K .......... .......... ........                        100%  213M=1.1s

2020-03-02 03:27:29 (6.97 Mb/s) - ‘/dev/null’ saved [951003/951003]

