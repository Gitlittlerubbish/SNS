--2020-02-25 22:12:32--  http://www.digestyc.gob.sv/EHPM2012/digestyc/resultado.pdf%0D
Resolving www.digestyc.gob.sv (www.digestyc.gob.sv)... 179.5.80.106
Connecting to www.digestyc.gob.sv (www.digestyc.gob.sv)|179.5.80.106|:80... failed: Connection timed out.
Giving up.

--2020-02-25 22:13:16--  http://www.digestyc.gob.sv/EHPM2012/digestyc/resultado.pdf%0D
Resolving www.digestyc.gob.sv (www.digestyc.gob.sv)... 179.5.80.106
Connecting to www.digestyc.gob.sv (www.digestyc.gob.sv)|179.5.80.106|:80... failed: Connection timed out.
Giving up.

