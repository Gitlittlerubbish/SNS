--2020-02-25 22:14:13--  http://www.ops.com.sv/pdf/205SESeries-Brochure.pdf%0D
Resolving www.ops.com.sv (www.ops.com.sv)... 192.185.148.211
Connecting to www.ops.com.sv (www.ops.com.sv)|192.185.148.211|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:14 ERROR 404: Not Found.

--2020-02-25 22:14:38--  http://www.ops.com.sv/pdf/205SESeries-Brochure.pdf%0D
Resolving www.ops.com.sv (www.ops.com.sv)... 192.185.148.211
Connecting to www.ops.com.sv (www.ops.com.sv)|192.185.148.211|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:38 ERROR 404: Not Found.

