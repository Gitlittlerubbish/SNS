--2020-02-25 22:14:00--  https://www.uees.edu.sv/carreras/pensumpdf/pensumnegociosinternacionales2.pdf%0D
Resolving www.uees.edu.sv (www.uees.edu.sv)... 201.162.197.198
Connecting to www.uees.edu.sv (www.uees.edu.sv)|201.162.197.198|:443... connected.
HTTP request sent, awaiting response... 404 Not found
2020-02-25 22:14:01 ERROR 404: Not found.

--2020-02-25 22:14:26--  https://www.uees.edu.sv/carreras/pensumpdf/pensumnegociosinternacionales2.pdf%0D
Resolving www.uees.edu.sv (www.uees.edu.sv)... 201.162.197.198
Connecting to www.uees.edu.sv (www.uees.edu.sv)|201.162.197.198|:443... connected.
HTTP request sent, awaiting response... 404 Not found
2020-02-25 22:14:28 ERROR 404: Not found.

