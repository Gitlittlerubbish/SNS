--2020-03-02 03:26:21--  http://santatecla.gob.sv/documentos/Servicios-Catastro.pdf
Resolving santatecla.gob.sv (santatecla.gob.sv)... 192.254.190.129
Connecting to santatecla.gob.sv (santatecla.gob.sv)|192.254.190.129|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 163050 (159K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 31% 1.20M 1s
    50K .......... .......... .......... .......... .......... 62% 2.44M 0s
   100K .......... .......... .......... .......... .......... 94% 67.6M 0s
   150K .........                                             100%  900M=0.5s

2020-03-02 03:26:23 (2.53 Mb/s) - ‘/dev/null’ saved [163050/163050]

