--2020-03-02 03:27:22--  http://www.qualitas.com.sv/web/qsv/red-talleres
Resolving www.qualitas.com.sv (www.qualitas.com.sv)... 190.86.175.251
Connecting to www.qualitas.com.sv (www.qualitas.com.sv)|190.86.175.251|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 336824 (329K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 15% 1.51M 2s
    50K .......... .......... .......... .......... .......... 30% 3.04M 1s
   100K .......... .......... .......... .......... .......... 45% 32.2M 0s
   150K .......... .......... .......... .......... .......... 60% 42.4M 0s
   200K .......... .......... .......... .......... .......... 76% 3.39M 0s
   250K .......... .......... .......... .......... .......... 91% 35.3M 0s
   300K .......... .......... ........                        100% 34.1M=0.6s

2020-03-02 03:27:26 (4.75 Mb/s) - ‘/dev/null’ saved [336824/336824]

