--2020-03-02 03:25:15--  http://www.cultura.gob.sv/wp-content/uploads/2016/08/Revista_ARS_10.pdf
Resolving www.cultura.gob.sv (www.cultura.gob.sv)... 190.120.4.18
Connecting to www.cultura.gob.sv (www.cultura.gob.sv)|190.120.4.18|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 15163002 (14M) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  0% 1.45M 83s
    50K .......... .......... .......... .......... ..........  0% 2.65M 64s
   100K .......... .......... .......... .......... ..........  1% 2.91M 56s
   150K .......... .......... .......... .......... ..........  1% 2.15M 56s
   200K .......... .......... .......... .......... ..........  1%  423M 45s
   250K .......... .......... .......... .......... ..........  2% 3.00M 44s
   300K .......... .......... .......... .......... ..........  2% 10.2M 39s
   350K .......... .......... .......... .......... ..........  2% 8.00M 36s
   400K .......... .......... .......... .......... ..........  3% 8.97M 33s
   450K .......... .......... .......... .......... ..........  3% 21.1M 30s
   500K .......... .......... .......... .......... ..........  3% 6.97M 29s
   550K .......... .......... .......... .......... ..........  4% 9.36M 28s
   600K .......... .......... .......... .......... ..........  4% 7.92M 26s
   650K .......... .......... .......... .......... ..........  4% 11.7M 25s
   700K .......... .......... .......... .......... ..........  5% 18.9M 24s
   750K .......... .......... .......... .......... ..........  5% 6.83M 23s
   800K .......... .......... .......... .......... ..........  5% 9.22M 23s
   850K .......... .......... .......... .......... ..........  6% 8.63M 22s
   900K .......... .......... .......... .......... ..........  6% 11.1M 21s
   950K .......... .......... .......... .......... ..........  6% 19.6M 20s
  1000K .......... .......... .......... .......... ..........  7% 6.80M 20s
  1050K .......... .......... .......... .......... ..........  7% 10.3M 20s
  1100K .......... .......... .......... .......... ..........  7% 10.4M 19s
  1150K .......... .......... .......... .......... ..........  8% 7.92M 19s
  1200K .......... .......... .......... .......... ..........  8% 20.4M 18s
  1250K .......... .......... .......... .......... ..........  8% 6.95M 18s
  1300K .......... .......... .......... .......... ..........  9% 9.11M 18s
  1350K .......... .......... .......... .......... ..........  9% 12.7M 18s
  1400K .......... .......... .......... .......... ..........  9% 11.9M 17s
  1450K .......... .......... .......... .......... .......... 10% 13.1M 17s
  1500K .......... .......... .......... .......... .......... 10% 6.95M 17s
  1550K .......... .......... .......... .......... .......... 10% 9.31M 16s
  1600K .......... .......... .......... .......... .......... 11% 8.89M 16s
  1650K .......... .......... .......... .......... .......... 11% 24.0M 16s
  1700K .......... .......... .......... .......... .......... 11% 9.99M 16s
  1750K .......... .......... .......... .......... .......... 12% 6.44M 16s
  1800K .......... .......... .......... .......... .......... 12% 9.84M 15s
  1850K .......... .......... .......... .......... .......... 12% 27.8M 15s
  1900K .......... .......... .......... .......... .......... 13% 9.53M 15s
  1950K .......... .......... .......... .......... .......... 13% 7.57M 15s
  2000K .......... .......... .......... .......... .......... 13% 7.08M 15s
  2050K .......... .......... .......... .......... .......... 14% 10.6M 15s
  2100K .......... .......... .......... .......... .......... 14% 22.0M 14s
  2150K .......... .......... .......... .......... .......... 14% 9.48M 14s
  2200K .......... .......... .......... .......... .......... 15% 6.39M 14s
  2250K .......... .......... .......... .......... .......... 15% 10.3M 14s
  2300K .......... .......... .......... .......... .......... 15% 8.63M 14s
  2350K .......... .......... .......... .......... .......... 16%  100M 14s
  2400K .......... .......... .......... .......... .......... 16% 5.93M 14s
  2450K .......... .......... .......... .......... .......... 16% 13.6M 13s
  2500K .......... .......... .......... .......... .......... 17% 8.69M 13s
  2550K .......... .......... .......... .......... .......... 17% 7.89M 13s
  2600K .......... .......... .......... .......... .......... 17%  160M 13s
  2650K .......... .......... .......... .......... .......... 18% 5.83M 13s
  2700K .......... .......... .......... .......... .......... 18% 9.79M 13s
  2750K .......... .......... .......... .......... .......... 18% 8.34M 13s
  2800K .......... .......... .......... .......... .......... 19% 9.59M 13s
  2850K .......... .......... .......... .......... .......... 19%  207M 12s
  2900K .......... .......... .......... .......... .......... 19% 6.55M 12s
  2950K .......... .......... .......... .......... .......... 20% 8.94M 12s
  3000K .......... .......... .......... .......... .......... 20% 8.10M 12s
  3050K .......... .......... .......... .......... .......... 20% 8.67M 12s
  3100K .......... .......... .......... .......... .......... 21%  144M 12s
  3150K .......... .......... .......... .......... .......... 21% 5.90M 12s
  3200K .......... .......... .......... .......... .......... 21% 9.73M 12s
  3250K .......... .......... .......... .......... .......... 22% 9.55M 12s
  3300K .......... .......... .......... .......... .......... 22% 7.94M 12s
  3350K .......... .......... .......... .......... .......... 22%  112M 12s
  3400K .......... .......... .......... .......... .......... 23% 5.26M 12s
  3450K .......... .......... .......... .......... .......... 23% 15.3M 12s
  3500K .......... .......... .......... .......... .......... 23% 7.84M 11s
  3550K .......... .......... .......... .......... .......... 24% 8.55M 11s
  3600K .......... .......... .......... .......... .......... 24%  133M 11s
  3650K .......... .......... .......... .......... .......... 24% 6.66M 11s
  3700K .......... .......... .......... .......... .......... 25% 9.43M 11s
  3750K .......... .......... .......... .......... .......... 25% 7.88M 11s
  3800K .......... .......... .......... .......... .......... 26% 8.03M 11s
  3850K .......... .......... .......... .......... .......... 26%  188M 11s
  3900K .......... .......... .......... .......... .......... 26% 6.08M 11s
  3950K .......... .......... .......... .......... .......... 27% 11.4M 11s
  4000K .......... .......... .......... .......... .......... 27% 7.76M 11s
  4050K .......... .......... .......... .......... .......... 27% 8.18M 11s
  4100K .......... .......... .......... .......... .......... 28% 40.9M 11s
  4150K .......... .......... .......... .......... .......... 28% 7.91M 10s
  4200K .......... .......... .......... .......... .......... 28% 9.31M 10s
  4250K .......... .......... .......... .......... .......... 29% 7.08M 10s
  4300K .......... .......... .......... .......... .......... 29% 9.13M 10s
  4350K .......... .......... .......... .......... .......... 29% 31.2M 10s
  4400K .......... .......... .......... .......... .......... 30% 7.27M 10s
  4450K .......... .......... .......... .......... .......... 30% 11.4M 10s
  4500K .......... .......... .......... .......... .......... 30% 4.51M 10s
  4550K .......... .......... .......... .......... .......... 31%  246M 10s
  4600K .......... .......... .......... .......... .......... 31% 8.03M 10s
  4650K .......... .......... .......... .......... .......... 31% 5.62M 10s
  4700K .......... .......... .......... .......... .......... 32% 13.6M 10s
  4750K .......... .......... .......... .......... .......... 32% 7.86M 10s
  4800K .......... .......... .......... .......... .......... 32%  207M 10s
  4850K .......... .......... .......... .......... .......... 33% 6.92M 10s
  4900K .......... .......... .......... .......... .......... 33% 5.93M 10s
  4950K .......... .......... .......... .......... .......... 33% 11.7M 10s
  5000K .......... .......... .......... .......... .......... 34% 9.60M 9s
  5050K .......... .......... .......... .......... .......... 34%  184M 9s
  5100K .......... .......... .......... .......... .......... 34% 6.59M 9s
  5150K .......... .......... .......... .......... .......... 35% 10.1M 9s
  5200K .......... .......... .......... .......... .......... 35% 6.33M 9s
  5250K .......... .......... .......... .......... .......... 35% 10.1M 9s
  5300K .......... .......... .......... .......... .......... 36%  236M 9s
  5350K .......... .......... .......... .......... .......... 36% 7.16M 9s
  5400K .......... .......... .......... .......... .......... 36% 9.31M 9s
  5450K .......... .......... .......... .......... .......... 37% 6.92M 9s
  5500K .......... .......... .......... .......... .......... 37% 9.33M 9s
  5550K .......... .......... .......... .......... .......... 37% 39.6M 9s
  5600K .......... .......... .......... .......... .......... 38% 8.85M 9s
  5650K .......... .......... .......... .......... .......... 38% 7.41M 9s
  5700K .......... .......... .......... .......... .......... 38% 7.13M 9s
  5750K .......... .......... .......... .......... .......... 39% 10.2M 9s
  5800K .......... .......... .......... .......... .......... 39% 34.6M 8s
  5850K .......... .......... .......... .......... .......... 39% 8.26M 8s
  5900K .......... .......... .......... .......... .......... 40% 9.63M 8s
  5950K .......... .......... .......... .......... .......... 40% 6.21M 8s
  6000K .......... .......... .......... .......... .......... 40% 10.5M 8s
  6050K .......... .......... .......... .......... .......... 41% 48.3M 8s
  6100K .......... .......... .......... .......... .......... 41% 8.76M 8s
  6150K .......... .......... .......... .......... .......... 41% 8.65M 8s
  6200K .......... .......... .......... .......... .......... 42% 6.69M 8s
  6250K .......... .......... .......... .......... .......... 42% 9.32M 8s
  6300K .......... .......... .......... .......... .......... 42% 24.5M 8s
  6350K .......... .......... .......... .......... .......... 43% 6.01M 8s
  6400K .......... .......... .......... .......... .......... 43% 22.6M 8s
  6450K .......... .......... .......... .......... .......... 43% 6.49M 8s
  6500K .......... .......... .......... .......... .......... 44% 10.3M 8s
  6550K .......... .......... .......... .......... .......... 44% 44.8M 8s
  6600K .......... .......... .......... .......... .......... 44% 7.41M 8s
  6650K .......... .......... .......... .......... .......... 45% 9.06M 8s
  6700K .......... .......... .......... .......... .......... 45% 8.39M 8s
  6750K .......... .......... .......... .......... .......... 45% 8.23M 7s
  6800K .......... .......... .......... .......... .......... 46% 90.3M 7s
  6850K .......... .......... .......... .......... .......... 46% 6.36M 7s
  6900K .......... .......... .......... .......... .......... 46% 11.0M 7s
  6950K .......... .......... .......... .......... .......... 47% 7.05M 7s
  7000K .......... .......... .......... .......... .......... 47% 9.32M 7s
  7050K .......... .......... .......... .......... .......... 47% 41.3M 7s
  7100K .......... .......... .......... .......... .......... 48% 6.46M 7s
  7150K .......... .......... .......... .......... .......... 48% 12.4M 7s
  7200K .......... .......... .......... .......... .......... 48% 6.58M 7s
  7250K .......... .......... .......... .......... .......... 49% 10.4M 7s
  7300K .......... .......... .......... .......... .......... 49%  129M 7s
  7350K .......... .......... .......... .......... .......... 49% 5.51M 7s
  7400K .......... .......... .......... .......... .......... 50% 11.5M 7s
  7450K .......... .......... .......... .......... .......... 50% 8.96M 7s
  7500K .......... .......... .......... .......... .......... 50% 6.71M 7s
  7550K .......... .......... .......... .......... .......... 51%  130M 7s
  7600K .......... .......... .......... .......... .......... 51% 5.61M 7s
  7650K .......... .......... .......... .......... .......... 52% 10.2M 7s
  7700K .......... .......... .......... .......... .......... 52% 8.67M 7s
  7750K .......... .......... .......... .......... .......... 52% 9.64M 6s
  7800K .......... .......... .......... .......... .......... 53% 30.5M 6s
  7850K .......... .......... .......... .......... .......... 53% 7.79M 6s
  7900K .......... .......... .......... .......... .......... 53% 7.04M 6s
  7950K .......... .......... .......... .......... .......... 54% 11.5M 6s
  8000K .......... .......... .......... .......... .......... 54%  121M 6s
  8050K .......... .......... .......... .......... .......... 54% 6.23M 6s
  8100K .......... .......... .......... .......... .......... 55% 11.1M 6s
  8150K .......... .......... .......... .......... .......... 55% 8.02M 6s
  8200K .......... .......... .......... .......... .......... 55% 8.09M 6s
  8250K .......... .......... .......... .......... .......... 56% 93.2M 6s
  8300K .......... .......... .......... .......... .......... 56% 7.06M 6s
  8350K .......... .......... .......... .......... .......... 56% 9.26M 6s
  8400K .......... .......... .......... .......... .......... 57% 7.93M 6s
  8450K .......... .......... .......... .......... .......... 57% 8.02M 6s
  8500K .......... .......... .......... .......... .......... 57% 9.43M 6s
  8550K .......... .......... .......... .......... .......... 58% 39.7M 6s
  8600K .......... .......... .......... .......... .......... 58% 7.94M 6s
  8650K .......... .......... .......... .......... .......... 58% 5.95M 6s
  8700K .......... .......... .......... .......... .......... 59% 12.2M 6s
  8750K .......... .......... .......... .......... .......... 59%  138M 5s
  8800K .......... .......... .......... .......... .......... 59% 8.03M 5s
  8850K .......... .......... .......... .......... .......... 60% 7.43M 5s
  8900K .......... .......... .......... .......... .......... 60% 8.64M 5s
  8950K .......... .......... .......... .......... .......... 60% 7.71M 5s
  9000K .......... .......... .......... .......... .......... 61% 1.23G 5s
  9050K .......... .......... .......... .......... .......... 61% 7.85M 5s
  9100K .......... .......... .......... .......... .......... 61% 7.99M 5s
  9150K .......... .......... .......... .......... .......... 62% 7.78M 5s
  9200K .......... .......... .......... .......... .......... 62% 8.01M 5s
  9250K .......... .......... .......... .......... .......... 62%  305M 5s
  9300K .......... .......... .......... .......... .......... 63% 7.41M 5s
  9350K .......... .......... .......... .......... .......... 63% 8.67M 5s
  9400K .......... .......... .......... .......... .......... 63% 7.86M 5s
  9450K .......... .......... .......... .......... .......... 64% 7.72M 5s
  9500K .......... .......... .......... .......... .......... 64% 39.4M 5s
  9550K .......... .......... .......... .......... .......... 64% 9.61M 5s
  9600K .......... .......... .......... .......... .......... 65% 8.19M 5s
  9650K .......... .......... .......... .......... .......... 65% 7.84M 5s
  9700K .......... .......... .......... .......... .......... 65% 8.11M 5s
  9750K .......... .......... .......... .......... .......... 66% 28.5M 5s
  9800K .......... .......... .......... .......... .......... 66% 9.27M 4s
  9850K .......... .......... .......... .......... .......... 66% 7.19M 4s
  9900K .......... .......... .......... .......... .......... 67% 7.96M 4s
  9950K .......... .......... .......... .......... .......... 67% 9.97M 4s
 10000K .......... .......... .......... .......... .......... 67% 22.9M 4s
 10050K .......... .......... .......... .......... .......... 68% 10.5M 4s
 10100K .......... .......... .......... .......... .......... 68% 6.53M 4s
 10150K .......... .......... .......... .......... .......... 68% 10.8M 4s
 10200K .......... .......... .......... .......... .......... 69% 8.07M 4s
 10250K .......... .......... .......... .......... .......... 69% 33.9M 4s
 10300K .......... .......... .......... .......... .......... 69% 8.14M 4s
 10350K .......... .......... .......... .......... .......... 70% 7.67M 4s
 10400K .......... .......... .......... .......... .......... 70% 9.96M 4s
 10450K .......... .......... .......... .......... .......... 70% 8.01M 4s
 10500K .......... .......... .......... .......... .......... 71% 9.71M 4s
 10550K .......... .......... .......... .......... .......... 71% 15.9M 4s
 10600K .......... .......... .......... .......... .......... 71% 7.42M 4s
 10650K .......... .......... .......... .......... .......... 72% 9.98M 4s
 10700K .......... .......... .......... .......... .......... 72% 9.19M 4s
 10750K .......... .......... .......... .......... .......... 72% 13.5M 4s
 10800K .......... .......... .......... .......... .......... 73% 9.19M 4s
 10850K .......... .......... .......... .......... .......... 73% 13.1M 3s
 10900K .......... .......... .......... .......... .......... 73% 8.02M 3s
 10950K .......... .......... .......... .......... .......... 74% 7.99M 3s
 11000K .......... .......... .......... .......... .......... 74% 10.2M 3s
 11050K .......... .......... .......... .......... .......... 74% 10.7M 3s
 11100K .......... .......... .......... .......... .......... 75% 11.5M 3s
 11150K .......... .......... .......... .......... .......... 75% 9.49M 3s
 11200K .......... .......... .......... .......... .......... 75% 9.69M 3s
 11250K .......... .......... .......... .......... .......... 76% 36.5M 3s
 11300K .......... .......... .......... .......... .......... 76% 5.21M 3s
 11350K .......... .......... .......... .......... .......... 76% 11.6M 3s
 11400K .......... .......... .......... .......... .......... 77% 10.3M 3s
 11450K .......... .......... .......... .......... .......... 77% 20.4M 3s
 11500K .......... .......... .......... .......... .......... 78% 9.86M 3s
 11550K .......... .......... .......... .......... .......... 78% 8.92M 3s
 11600K .......... .......... .......... .......... .......... 78% 6.73M 3s
 11650K .......... .......... .......... .......... .......... 79% 10.0M 3s
 11700K .......... .......... .......... .......... .......... 79% 17.8M 3s
 11750K .......... .......... .......... .......... .......... 79% 13.2M 3s
 11800K .......... .......... .......... .......... .......... 80% 8.17M 3s
 11850K .......... .......... .......... .......... .......... 80% 6.14M 3s
 11900K .......... .......... .......... .......... .......... 80% 11.1M 3s
 11950K .......... .......... .......... .......... .......... 81% 15.5M 2s
 12000K .......... .......... .......... .......... .......... 81% 12.0M 2s
 12050K .......... .......... .......... .......... .......... 81% 9.22M 2s
 12100K .......... .......... .......... .......... .......... 82% 7.95M 2s
 12150K .......... .......... .......... .......... .......... 82% 7.89M 2s
 12200K .......... .......... .......... .......... .......... 82% 26.4M 2s
 12250K .......... .......... .......... .......... .......... 83% 8.30M 2s
 12300K .......... .......... .......... .......... .......... 83% 10.2M 2s
 12350K .......... .......... .......... .......... .......... 83% 8.07M 2s
 12400K .......... .......... .......... .......... .......... 84% 7.67M 2s
 12450K .......... .......... .......... .......... .......... 84% 44.1M 2s
 12500K .......... .......... .......... .......... .......... 84% 7.09M 2s
 12550K .......... .......... .......... .......... .......... 85% 11.4M 2s
 12600K .......... .......... .......... .......... .......... 85% 7.87M 2s
 12650K .......... .......... .......... .......... .......... 85% 8.07M 2s
 12700K .......... .......... .......... .......... .......... 86% 21.3M 2s
 12750K .......... .......... .......... .......... .......... 86% 9.47M 2s
 12800K .......... .......... .......... .......... .......... 86% 9.46M 2s
 12850K .......... .......... .......... .......... .......... 87% 6.84M 2s
 12900K .......... .......... .......... .......... .......... 87% 9.56M 2s
 12950K .......... .......... .......... .......... .......... 87% 16.7M 2s
 13000K .......... .......... .......... .......... .......... 88% 10.0M 2s
 13050K .......... .......... .......... .......... .......... 88% 10.2M 2s
 13100K .......... .......... .......... .......... .......... 88% 8.00M 1s
 13150K .......... .......... .......... .......... .......... 89% 7.89M 1s
 13200K .......... .......... .......... .......... .......... 89% 18.6M 1s
 13250K .......... .......... .......... .......... .......... 89% 10.3M 1s
 13300K .......... .......... .......... .......... .......... 90% 9.40M 1s
 13350K .......... .......... .......... .......... .......... 90% 7.94M 1s
 13400K .......... .......... .......... .......... .......... 90% 8.11M 1s
 13450K .......... .......... .......... .......... .......... 91% 5.09M 1s
 13500K .......... .......... .......... .......... .......... 91%  155M 1s
 13550K .......... .......... .......... .......... .......... 91% 13.1M 1s
 13600K .......... .......... .......... .......... .......... 92% 8.10M 1s
 13650K .......... .......... .......... .......... .......... 92% 9.34M 1s
 13700K .......... .......... .......... .......... .......... 92% 32.7M 1s
 13750K .......... .......... .......... .......... .......... 93% 9.50M 1s
 13800K .......... .......... .......... .......... .......... 93% 8.07M 1s
 13850K .......... .......... .......... .......... .......... 93% 7.99M 1s
 13900K .......... .......... .......... .......... .......... 94% 8.04M 1s
 13950K .......... .......... .......... .......... .......... 94%  139M 1s
 14000K .......... .......... .......... .......... .......... 94% 7.05M 1s
 14050K .......... .......... .......... .......... .......... 95% 8.34M 1s
 14100K .......... .......... .......... .......... .......... 95% 7.64M 1s
 14150K .......... .......... .......... .......... .......... 95% 9.34M 1s
 14200K .......... .......... .......... .......... .......... 96%  104M 0s
 14250K .......... .......... .......... .......... .......... 96% 8.23M 0s
 14300K .......... .......... .......... .......... .......... 96% 7.74M 0s
 14350K .......... .......... .......... .......... .......... 97% 8.13M 0s
 14400K .......... .......... .......... .......... .......... 97%  193M 0s
 14450K .......... .......... .......... .......... .......... 97% 6.51M 0s
 14500K .......... .......... .......... .......... .......... 98% 8.11M 0s
 14550K .......... .......... .......... .......... .......... 98% 9.73M 0s
 14600K .......... .......... .......... .......... .......... 98% 7.93M 0s
 14650K .......... .......... .......... .......... .......... 99% 34.6M 0s
 14700K .......... .......... .......... .......... .......... 99% 7.29M 0s
 14750K .......... .......... .......... .......... .......... 99% 9.07M 0s
 14800K .......                                               100% 2.48M=13s

2020-03-02 03:25:31 (9.32 Mb/s) - ‘/dev/null’ saved [15163002/15163002]

