--2020-02-25 22:13:43--  http://www.minsal.sv/archivos/chagas2008/pdf/La_enfermedad_de_chagas_en_el_salvador_evolucion_historica_y_desafio_para_el_control.pdf%0D
Resolving www.minsal.sv (www.minsal.sv)... 190.86.223.123
Connecting to www.minsal.sv (www.minsal.sv)|190.86.223.123|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:45 ERROR 404: Not Found.

--2020-02-25 22:14:13--  http://www.minsal.sv/archivos/chagas2008/pdf/La_enfermedad_de_chagas_en_el_salvador_evolucion_historica_y_desafio_para_el_control.pdf%0D
Resolving www.minsal.sv (www.minsal.sv)... 190.86.223.123
Connecting to www.minsal.sv (www.minsal.sv)|190.86.223.123|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:15 ERROR 404: Not Found.

