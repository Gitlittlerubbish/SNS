--2020-03-02 03:24:17--  http://tramites.gob.sv/media/Codigo_municipal.pdf
Resolving tramites.gob.sv (tramites.gob.sv)... 136.243.24.150
Connecting to tramites.gob.sv (tramites.gob.sv)|136.243.24.150|:80... connected.
HTTP request sent, awaiting response... 302 Redirect
Location: https://tramites.gob.sv/media/Codigo_municipal.pdf [following]
--2020-03-02 03:24:17--  https://tramites.gob.sv/media/Codigo_municipal.pdf
Connecting to tramites.gob.sv (tramites.gob.sv)|136.243.24.150|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: 243466 (238K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 21% 9.39M 0s
    50K .......... .......... .......... .......... .......... 42% 84.2M 0s
   100K .......... .......... .......... .......... .......... 63% 17.8M 0s
   150K .......... .......... .......... .......... .......... 84%  196M 0s
   200K .......... .......... .......... .......              100%  275M=0.07s

2020-03-02 03:24:17 (26.1 Mb/s) - ‘/dev/null’ saved [243466/243466]

