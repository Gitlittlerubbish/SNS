--2020-03-02 03:23:58--  http://www.yamaha-motor.com.sv/home/storage/documents/QvbsNSQyqeaYdfIBTUK5KxEZCJEDABeZlmzDjQXM.pdf
Resolving www.yamaha-motor.com.sv (www.yamaha-motor.com.sv)... 72.47.228.69
Connecting to www.yamaha-motor.com.sv (www.yamaha-motor.com.sv)|72.47.228.69|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 4542489 (4.3M) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  1% 1.45M 25s
    50K .......... .......... .......... .......... ..........  2% 2.93M 18s
   100K .......... .......... .......... .......... ..........  3%  110M 12s
   150K .......... .......... .......... .......... ..........  4%  146M 9s
   200K .......... .......... .......... .......... ..........  5% 2.94M 10s
   250K .......... .......... .......... .......... ..........  6%  180M 8s
   300K .......... .......... .......... .......... ..........  7% 2.92M 8s
   350K .......... .......... .......... .......... ..........  9%  141M 7s
   400K .......... .......... .......... .......... .......... 10%  531M 6s
   450K .......... .......... .......... .......... .......... 11%  340M 6s
   500K .......... .......... .......... .......... .......... 12%  133M 5s
   550K .......... .......... .......... .......... .......... 13% 3.06M 5s
   600K .......... .......... .......... .......... .......... 14% 83.3M 5s
   650K .......... .......... .......... .......... .......... 15%  164M 5s
   700K .......... .......... .......... .......... .......... 16%  407M 4s
   750K .......... .......... .......... .......... .......... 18%  314M 4s
   800K .......... .......... .......... .......... .......... 19% 3.10M 4s
   850K .......... .......... .......... .......... .......... 20%  214M 4s
   900K .......... .......... .......... .......... .......... 21%  350M 4s
   950K .......... .......... .......... .......... .......... 22%  277M 3s
  1000K .......... .......... .......... .......... .......... 23%  304M 3s
  1050K .......... .......... .......... .......... .......... 24%  107M 3s
  1100K .......... .......... .......... .......... .......... 25%  483M 3s
  1150K .......... .......... .......... .......... .......... 27% 4.09M 3s
  1200K .......... .......... .......... .......... .......... 28% 14.6M 3s
  1250K .......... .......... .......... .......... .......... 29%  212M 3s
  1300K .......... .......... .......... .......... .......... 30% 66.7M 3s
  1350K .......... .......... .......... .......... .......... 31%  363M 2s
  1400K .......... .......... .......... .......... .......... 32%  262M 2s
  1450K .......... .......... .......... .......... .......... 33%  184M 2s
  1500K .......... .......... .......... .......... .......... 34%  230M 2s
  1550K .......... .......... .......... .......... .......... 36%  200M 2s
  1600K .......... .......... .......... .......... .......... 37%  488M 2s
  1650K .......... .......... .......... .......... .......... 38% 3.26M 2s
  1700K .......... .......... .......... .......... .......... 39%  232M 2s
  1750K .......... .......... .......... .......... .......... 40%  274M 2s
  1800K .......... .......... .......... .......... .......... 41%  139M 2s
  1850K .......... .......... .......... .......... .......... 42%  588M 2s
  1900K .......... .......... .......... .......... .......... 43%  219M 2s
  1950K .......... .......... .......... .......... .......... 45%  159M 2s
  2000K .......... .......... .......... .......... .......... 46% 1.08G 1s
  2050K .......... .......... .......... .......... .......... 47%  182M 1s
  2100K .......... .......... .......... .......... .......... 48%  587M 1s
  2150K .......... .......... .......... .......... .......... 49%  213M 1s
  2200K .......... .......... .......... .......... .......... 50%  374M 1s
  2250K .......... .......... .......... .......... .......... 51%  277M 1s
  2300K .......... .......... .......... .......... .......... 52%  210M 1s
  2350K .......... .......... .......... .......... .......... 54%  455M 1s
  2400K .......... .......... .......... .......... .......... 55%  385M 1s
  2450K .......... .......... .......... .......... .......... 56%  121M 1s
  2500K .......... .......... .......... .......... .......... 57% 3.28M 1s
  2550K .......... .......... .......... .......... .......... 58%  528M 1s
  2600K .......... .......... .......... .......... .......... 59%  249M 1s
  2650K .......... .......... .......... .......... .......... 60%  339M 1s
  2700K .......... .......... .......... .......... .......... 61%  335M 1s
  2750K .......... .......... .......... .......... .......... 63%  231M 1s
  2800K .......... .......... .......... .......... .......... 64%  198M 1s
  2850K .......... .......... .......... .......... .......... 65%  356M 1s
  2900K .......... .......... .......... .......... .......... 66%  361M 1s
  2950K .......... .......... .......... .......... .......... 67%  260M 1s
  3000K .......... .......... .......... .......... .......... 68%  390M 1s
  3050K .......... .......... .......... .......... .......... 69%  188M 1s
  3100K .......... .......... .......... .......... .......... 71%  256M 1s
  3150K .......... .......... .......... .......... .......... 72%  329M 1s
  3200K .......... .......... .......... .......... .......... 73%  429M 1s
  3250K .......... .......... .......... .......... .......... 74%  217M 0s
  3300K .......... .......... .......... .......... .......... 75%  565M 0s
  3350K .......... .......... .......... .......... .......... 76%  191M 0s
  3400K .......... .......... .......... .......... .......... 77%  331M 0s
  3450K .......... .......... .......... .......... .......... 78% 3.70M 0s
  3500K .......... .......... .......... .......... .......... 80% 38.5M 0s
  3550K .......... .......... .......... .......... .......... 81%  159M 0s
  3600K .......... .......... .......... .......... .......... 82%  206M 0s
  3650K .......... .......... .......... .......... .......... 83%  467M 0s
  3700K .......... .......... .......... .......... .......... 84%  441M 0s
  3750K .......... .......... .......... .......... .......... 85%  405M 0s
  3800K .......... .......... .......... .......... .......... 86%  178M 0s
  3850K .......... .......... .......... .......... .......... 87%  210M 0s
  3900K .......... .......... .......... .......... .......... 89%  492M 0s
  3950K .......... .......... .......... .......... .......... 90%  464M 0s
  4000K .......... .......... .......... .......... .......... 91%  292M 0s
  4050K .......... .......... .......... .......... .......... 92%  107M 0s
  4100K .......... .......... .......... .......... .......... 93%  261M 0s
  4150K .......... .......... .......... .......... .......... 94% 2.80M 0s
  4200K .......... .......... .......... .......... .......... 95% 1.49G 0s
  4250K .......... .......... .......... .......... .......... 96% 1.32G 0s
  4300K .......... .......... .......... .......... .......... 98% 1.85G 0s
  4350K .......... .......... .......... .......... .......... 99% 1.88G 0s
  4400K .......... .......... .......... ......               100% 1.72G=1.7s

2020-03-02 03:24:01 (20.9 Mb/s) - ‘/dev/null’ saved [4542489/4542489]

