--2020-02-25 22:12:24--  http://www.psicopedagogico.edu.sv/archivoL/Libro009.pdf%0D
Resolving www.psicopedagogico.edu.sv (www.psicopedagogico.edu.sv)... failed: Connection timed out.
wget: unable to resolve host address ‘www.psicopedagogico.edu.sv’
--2020-02-25 22:13:14--  http://www.psicopedagogico.edu.sv/archivoL/Libro009.pdf%0D
Resolving www.psicopedagogico.edu.sv (www.psicopedagogico.edu.sv)... 66.7.198.130
Connecting to www.psicopedagogico.edu.sv (www.psicopedagogico.edu.sv)|66.7.198.130|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:15 ERROR 404: Not Found.

