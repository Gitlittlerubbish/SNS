--2020-03-02 03:23:53--  http://www.uca.edu.sv/-pDIq89
Resolving www.uca.edu.sv (www.uca.edu.sv)... 201.131.110.4
Connecting to www.uca.edu.sv (www.uca.edu.sv)|201.131.110.4|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 290 [text/html]
Saving to: ‘/dev/null’

     0K                                                       100%  116M=0s

2020-03-02 03:23:54 (116 Mb/s) - ‘/dev/null’ saved [290/290]

--2020-03-02 03:23:54--  http://www.uca.edu.sv/-1DUgTd
Resolving www.uca.edu.sv (www.uca.edu.sv)... 201.131.110.4
Connecting to www.uca.edu.sv (www.uca.edu.sv)|201.131.110.4|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 274 [text/html]
Saving to: ‘/dev/null’

     0K                                                       100% 78.3M=0s

2020-03-02 03:23:54 (78.3 Mb/s) - ‘/dev/null’ saved [274/274]

