--2020-02-25 22:12:49--  http://richmond.com.sv/ss/SSpathwaytoscience_g.pdf%0D
Resolving richmond.com.sv (richmond.com.sv)... 34.225.172.62, 34.238.101.91
Connecting to richmond.com.sv (richmond.com.sv)|34.225.172.62|:80... connected.
HTTP request sent, awaiting response... 404 Category not found
2020-02-25 22:12:50 ERROR 404: Category not found.

--2020-02-25 22:13:27--  http://richmond.com.sv/ss/SSpathwaytoscience_g.pdf%0D
Resolving richmond.com.sv (richmond.com.sv)... 34.225.172.62, 34.238.101.91
Connecting to richmond.com.sv (richmond.com.sv)|34.225.172.62|:80... connected.
HTTP request sent, awaiting response... 404 Category not found
2020-02-25 22:13:27 ERROR 404: Category not found.

