--2020-02-25 22:12:52--  https://tramites.gob.sv/media/Codigo_municipal.pdf%0D
Resolving tramites.gob.sv (tramites.gob.sv)... 136.243.24.150
Connecting to tramites.gob.sv (tramites.gob.sv)|136.243.24.150|:443... connected.
HTTP request sent, awaiting response... 400 Bad Request
2020-02-25 22:12:52 ERROR 400: Bad Request.

--2020-02-25 22:13:28--  https://tramites.gob.sv/media/Codigo_municipal.pdf%0D
Resolving tramites.gob.sv (tramites.gob.sv)... 136.243.24.150
Connecting to tramites.gob.sv (tramites.gob.sv)|136.243.24.150|:443... connected.
HTTP request sent, awaiting response... 400 Bad Request
2020-02-25 22:13:28 ERROR 400: Bad Request.

