--2020-03-02 03:27:20--  http://www.comures.org.sv/CIRCULAR-043-2017.pdf
Resolving www.comures.org.sv (www.comures.org.sv)... 174.142.89.94
Connecting to www.comures.org.sv (www.comures.org.sv)|174.142.89.94|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 255007 (249K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 20% 2.22M 1s
    50K .......... .......... .......... .......... .......... 40% 4.44M 0s
   100K .......... .......... .......... .......... .......... 60% 62.6M 0s
   150K .......... .......... .......... .......... .......... 80% 4.48M 0s
   200K .......... .......... .......... .......... ......... 100% 4.62M=0.5s

2020-03-02 03:27:22 (4.42 Mb/s) - ‘/dev/null’ saved [255007/255007]

