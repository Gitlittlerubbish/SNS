--2020-02-25 22:12:50--  http://www.amway.com.sv/downloads/Catalogo_Nutrilite_2015.pdf%0D
Resolving www.amway.com.sv (www.amway.com.sv)... 104.103.177.15
Connecting to www.amway.com.sv (www.amway.com.sv)|104.103.177.15|:80... connected.
HTTP request sent, awaiting response... 400 Bad Request
2020-02-25 22:12:51 ERROR 400: Bad Request.

--2020-02-25 22:13:27--  http://www.amway.com.sv/downloads/Catalogo_Nutrilite_2015.pdf%0D
Resolving www.amway.com.sv (www.amway.com.sv)... 104.103.177.15
Connecting to www.amway.com.sv (www.amway.com.sv)|104.103.177.15|:80... connected.
HTTP request sent, awaiting response... 400 Bad Request
2020-02-25 22:13:28 ERROR 400: Bad Request.

