--2020-03-02 03:23:54--  http://www.ufg.edu.sv/doc/FT-EBSCOhost.pdf
Resolving www.ufg.edu.sv (www.ufg.edu.sv)... 200.124.138.25
Connecting to www.ufg.edu.sv (www.ufg.edu.sv)|200.124.138.25|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 99488 (97K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 51% 1.47M 0s
    50K .......... .......... .......... .......... .......   100% 1.40M=0.6s

2020-03-02 03:23:56 (1.43 Mb/s) - ‘/dev/null’ saved [99488/99488]

