--2020-03-02 03:24:59--  http://www.upan.edu.sv/pdf/catalogo2017.pdf
Resolving www.upan.edu.sv (www.upan.edu.sv)... 143.95.150.52
Connecting to www.upan.edu.sv (www.upan.edu.sv)|143.95.150.52|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 2029149 (1.9M) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  2%  837K 19s
    50K .......... .......... .......... .......... ..........  5%  656K 21s
   100K .......... .......... .......... .......... ..........  7% 3.21M 15s
   150K .......... .......... .......... .......... .......... 10% 3.25M 12s
   200K .......... .......... .......... .......... .......... 12% 3.72M 10s
   250K .......... .......... .......... .......... .......... 15%  765K 11s
   300K .......... .......... .......... .......... .......... 17%  260M 9s
   350K .......... .......... .......... .......... .......... 20%  139M 8s
   400K .......... .......... .......... .......... .......... 22% 2.00M 8s
   450K .......... .......... .......... .......... .......... 25% 2.04M 7s
   500K .......... .......... .......... .......... .......... 27%  351M 6s
   550K .......... .......... .......... .......... .......... 30% 3.50M 6s
   600K .......... .......... .......... .......... .......... 32% 51.8M 5s
   650K .......... .......... .......... .......... .......... 35%  693K 6s
   700K .......... .......... .......... .......... .......... 37%  514M 5s
   750K .......... .......... .......... .......... .......... 40%  414M 5s
   800K .......... .......... .......... .......... .......... 42%  361M 4s
   850K .......... .......... .......... .......... .......... 45% 2.01M 4s
   900K .......... .......... .......... .......... .......... 47%  241M 4s
   950K .......... .......... .......... .......... .......... 50%  245M 3s
  1000K .......... .......... .......... .......... .......... 52% 2.04M 3s
  1050K .......... .......... .......... .......... .......... 55%  235M 3s
  1100K .......... .......... .......... .......... .......... 58%  389M 3s
  1150K .......... .......... .......... .......... .......... 60%  375M 2s
  1200K .......... .......... .......... .......... .......... 63%  167M 2s
  1250K .......... .......... .......... .......... .......... 65%  363M 2s
  1300K .......... .......... .......... .......... .......... 68% 3.42M 2s
  1350K .......... .......... .......... .......... .......... 70% 77.5M 2s
  1400K .......... .......... .......... .......... .......... 73%  101M 1s
  1450K .......... .......... .......... .......... .......... 75% 71.5M 1s
  1500K .......... .......... .......... .......... .......... 78% 59.0M 1s
  1550K .......... .......... .......... .......... .......... 80%  164M 1s
  1600K .......... .......... .......... .......... .......... 83% 5.10M 1s
  1650K .......... .......... .......... .......... .......... 85% 50.1M 1s
  1700K .......... .......... .......... .......... .......... 88% 82.5M 1s
  1750K .......... .......... .......... .......... .......... 90%  174M 0s
  1800K .......... .......... .......... .......... .......... 93%  154M 0s
  1850K .......... .......... .......... .......... .......... 95% 42.4M 0s
  1900K .......... .......... .......... .......... .......... 98%  103M 0s
  1950K .......... .......... .......... .                    100% 92.9M=3.8s

2020-03-02 03:25:04 (4.25 Mb/s) - ‘/dev/null’ saved [2029149/2029149]

