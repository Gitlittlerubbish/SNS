--2020-03-02 03:26:06--  http://www.cnr.gob.sv/documentos/igcn/requisitos_y_aranceles_de_servicio_.pdf
Resolving www.cnr.gob.sv (www.cnr.gob.sv)... 138.97.141.23
Connecting to www.cnr.gob.sv (www.cnr.gob.sv)|138.97.141.23|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: https://www.cnr.gob.sv/documentos/igcn/requisitos_y_aranceles_de_servicio_.pdf [following]
--2020-03-02 03:26:06--  https://www.cnr.gob.sv/documentos/igcn/requisitos_y_aranceles_de_servicio_.pdf
Connecting to www.cnr.gob.sv (www.cnr.gob.sv)|138.97.141.23|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: 797853 (779K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  6% 1.48M 4s
    50K .......... .......... .......... .......... .......... 12% 2.99M 3s
   100K .......... .......... .......... .......... .......... 19%  107M 2s
   150K .......... .......... .......... .......... .......... 25% 3.06M 2s
   200K .......... .......... .......... .......... .......... 32%  127M 1s
   250K .......... .......... .......... .......... .......... 38% 3.10M 1s
   300K .......... .......... .......... .......... .......... 44%  216M 1s
   350K .......... .......... .......... .......... .......... 51%  164M 1s
   400K .......... .......... .......... .......... .......... 57% 3.14M 1s
   450K .......... .......... .......... .......... .......... 64%  115M 0s
   500K .......... .......... .......... .......... .......... 70%  150M 0s
   550K .......... .......... .......... .......... .......... 77%  179M 0s
   600K .......... .......... .......... .......... .......... 83%  191M 0s
   650K .......... .......... .......... .......... .......... 89% 3.14M 0s
   700K .......... .......... .......... .......... .......... 96%  131M 0s
   750K .......... .......... .........                       100%  370M=1.0s

2020-03-02 03:26:08 (6.61 Mb/s) - ‘/dev/null’ saved [797853/797853]

