--2020-02-25 22:14:15--  http://www.qualitas.com.sv/web/qsv/red-talleres%0D
Resolving www.qualitas.com.sv (www.qualitas.com.sv)... 190.86.175.251
Connecting to www.qualitas.com.sv (www.qualitas.com.sv)|190.86.175.251|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:18 ERROR 404: Not Found.

--2020-02-25 22:14:39--  http://www.qualitas.com.sv/web/qsv/red-talleres%0D
Resolving www.qualitas.com.sv (www.qualitas.com.sv)... 190.86.175.251
Connecting to www.qualitas.com.sv (www.qualitas.com.sv)|190.86.175.251|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:39 ERROR 404: Not Found.

