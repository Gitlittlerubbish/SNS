--2020-03-02 03:25:31--  http://aplicaciones.itca.edu.sv/PwdCorreoITCA.pdf
Resolving aplicaciones.itca.edu.sv (aplicaciones.itca.edu.sv)... 200.35.188.115
Connecting to aplicaciones.itca.edu.sv (aplicaciones.itca.edu.sv)|200.35.188.115|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 788554 (770K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  6% 1.53M 4s
    50K .......... .......... .......... .......... .......... 12% 2.99M 3s
   100K .......... .......... .......... .......... .......... 19% 3.04M 2s
   150K .......... .......... .......... .......... .......... 25% 1.50M 2s
   200K .......... .......... .......... .......... .......... 32% 1.04G 2s
   250K .......... .......... .......... .......... .......... 38% 1.02M 2s
   300K .......... .......... .......... .......... .......... 45% 1.51M 2s
   350K .......... .......... .......... .......... .......... 51% 1.55M 2s
   400K .......... .......... .......... .......... .......... 58% 62.2M 1s
   450K .......... .......... .......... .......... .......... 64% 2.95M 1s
   500K .......... .......... .......... .......... .......... 71% 3.29M 1s
   550K .......... .......... .......... .......... .......... 77% 27.0M 1s
   600K .......... .......... .......... .......... .......... 84% 1.62M 0s
   650K .......... .......... .......... .......... .......... 90% 21.6M 0s
   700K .......... .......... .......... .......... .......... 97% 1.61M 0s
   750K .......... ..........                                 100% 13.2M=2.6s

2020-03-02 03:25:35 (2.45 Mb/s) - ‘/dev/null’ saved [788554/788554]

