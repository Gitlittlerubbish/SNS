--2020-02-25 22:14:20--  http://www.uma.edu.sv/image/pdf/diplomado.pdf%0D
Resolving www.uma.edu.sv (www.uma.edu.sv)... 200.30.138.51
Connecting to www.uma.edu.sv (www.uma.edu.sv)|200.30.138.51|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:21 ERROR 404: Not Found.

--2020-02-25 22:14:40--  http://www.uma.edu.sv/image/pdf/diplomado.pdf%0D
Resolving www.uma.edu.sv (www.uma.edu.sv)... 200.30.138.51
Connecting to www.uma.edu.sv (www.uma.edu.sv)|200.30.138.51|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:40 ERROR 404: Not Found.

