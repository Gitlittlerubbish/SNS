--2020-02-25 22:13:42--  http://www.evivienda.gob.sv/Lotificaciones/Documentos/INSTRUCTIVO_SIL.pdf%0D
Resolving www.evivienda.gob.sv (www.evivienda.gob.sv)... 200.31.181.149
Connecting to www.evivienda.gob.sv (www.evivienda.gob.sv)|200.31.181.149|:80... connected.
HTTP request sent, awaiting response... 400 Bad Request
2020-02-25 22:13:43 ERROR 400: Bad Request.

--2020-02-25 22:14:11--  http://www.evivienda.gob.sv/Lotificaciones/Documentos/INSTRUCTIVO_SIL.pdf%0D
Resolving www.evivienda.gob.sv (www.evivienda.gob.sv)... 200.31.181.149
Connecting to www.evivienda.gob.sv (www.evivienda.gob.sv)|200.31.181.149|:80... connected.
HTTP request sent, awaiting response... 400 Bad Request
2020-02-25 22:14:13 ERROR 400: Bad Request.

