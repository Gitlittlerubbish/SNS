--2020-03-02 03:24:05--  http://www.alges.org.sv/asset/documents/555
Resolving www.alges.org.sv (www.alges.org.sv)... 46.4.127.171
Connecting to www.alges.org.sv (www.alges.org.sv)|46.4.127.171|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... ..........                       10.1M=0.02s

2020-03-02 03:24:05 (10.1 Mb/s) - ‘/dev/null’ saved [30726]

