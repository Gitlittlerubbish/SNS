--2020-02-25 22:12:45--  http://www.innovacion.gob.sv/inventa/attachments/article/3569/cqb051e.pdf%0D
Resolving www.innovacion.gob.sv (www.innovacion.gob.sv)... 190.120.4.4
Connecting to www.innovacion.gob.sv (www.innovacion.gob.sv)|190.120.4.4|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: https://www.innovacion.gob.sv/inventa/attachments/article/3569/cqb051e.pdf%0d [following]
--2020-02-25 22:12:46--  https://www.innovacion.gob.sv/inventa/attachments/article/3569/cqb051e.pdf%0d
Connecting to www.innovacion.gob.sv (www.innovacion.gob.sv)|190.120.4.4|:443... connected.
ERROR: cannot verify www.innovacion.gob.sv's certificate, issued by ‘CN=Go Daddy Secure Certificate Authority - G2,OU=http://certs.godaddy.com/repository/,O=GoDaddy.com\\, Inc.,L=Scottsdale,ST=Arizona,C=US’:
  Unable to locally verify the issuer's authority.
To connect to www.innovacion.gob.sv insecurely, use `--no-check-certificate'.
--2020-02-25 22:13:24--  http://www.innovacion.gob.sv/inventa/attachments/article/3569/cqb051e.pdf%0D
Resolving www.innovacion.gob.sv (www.innovacion.gob.sv)... 190.120.4.4
Connecting to www.innovacion.gob.sv (www.innovacion.gob.sv)|190.120.4.4|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: https://www.innovacion.gob.sv/inventa/attachments/article/3569/cqb051e.pdf%0d [following]
--2020-02-25 22:13:24--  https://www.innovacion.gob.sv/inventa/attachments/article/3569/cqb051e.pdf%0d
Connecting to www.innovacion.gob.sv (www.innovacion.gob.sv)|190.120.4.4|:443... connected.
ERROR: cannot verify www.innovacion.gob.sv's certificate, issued by ‘CN=Go Daddy Secure Certificate Authority - G2,OU=http://certs.godaddy.com/repository/,O=GoDaddy.com\\, Inc.,L=Scottsdale,ST=Arizona,C=US’:
  Unable to locally verify the issuer's authority.
To connect to www.innovacion.gob.sv insecurely, use `--no-check-certificate'.
