--2020-02-25 22:13:50--  https://biblioteca.rree.gob.sv/textocompleto/271.pdf%0D
Resolving biblioteca.rree.gob.sv (biblioteca.rree.gob.sv)... 168.243.204.25
Connecting to biblioteca.rree.gob.sv (biblioteca.rree.gob.sv)|168.243.204.25|:443... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:53 ERROR 404: Not Found.

--2020-02-25 22:14:19--  https://biblioteca.rree.gob.sv/textocompleto/271.pdf%0D
Resolving biblioteca.rree.gob.sv (biblioteca.rree.gob.sv)... 168.243.204.25
Connecting to biblioteca.rree.gob.sv (biblioteca.rree.gob.sv)|168.243.204.25|:443... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:20 ERROR 404: Not Found.

