--2020-02-25 22:13:48--  http://www.cnr.gob.sv/documentos/igcn/requisitos_y_aranceles_de_servicio_.pdf%0D
Resolving www.cnr.gob.sv (www.cnr.gob.sv)... 138.97.141.23
Connecting to www.cnr.gob.sv (www.cnr.gob.sv)|138.97.141.23|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: https://www.cnr.gob.sv/documentos/igcn/requisitos_y_aranceles_de_servicio_.pdf%0d [following]
--2020-02-25 22:13:48--  https://www.cnr.gob.sv/documentos/igcn/requisitos_y_aranceles_de_servicio_.pdf%0d
Connecting to www.cnr.gob.sv (www.cnr.gob.sv)|138.97.141.23|:443... connected.
HTTP request sent, awaiting response... 403 Forbidden
2020-02-25 22:13:49 ERROR 403: Forbidden.

--2020-02-25 22:14:18--  http://www.cnr.gob.sv/documentos/igcn/requisitos_y_aranceles_de_servicio_.pdf%0D
Resolving www.cnr.gob.sv (www.cnr.gob.sv)... 138.97.141.23
Connecting to www.cnr.gob.sv (www.cnr.gob.sv)|138.97.141.23|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: https://www.cnr.gob.sv/documentos/igcn/requisitos_y_aranceles_de_servicio_.pdf%0d [following]
--2020-02-25 22:14:18--  https://www.cnr.gob.sv/documentos/igcn/requisitos_y_aranceles_de_servicio_.pdf%0d
Connecting to www.cnr.gob.sv (www.cnr.gob.sv)|138.97.141.23|:443... connected.
HTTP request sent, awaiting response... 403 Forbidden
2020-02-25 22:14:19 ERROR 403: Forbidden.

