--2020-02-25 22:14:19--  http://www.csj.gob.sv/INV_PROF/INV_PROF/TRAMITE_AA_22_11_12.pdf%0D
Resolving www.csj.gob.sv (www.csj.gob.sv)... 200.31.169.70
Connecting to www.csj.gob.sv (www.csj.gob.sv)|200.31.169.70|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:20 ERROR 404: Not Found.

--2020-02-25 22:14:39--  http://www.csj.gob.sv/INV_PROF/INV_PROF/TRAMITE_AA_22_11_12.pdf%0D
Resolving www.csj.gob.sv (www.csj.gob.sv)... 200.31.169.70
Connecting to www.csj.gob.sv (www.csj.gob.sv)|200.31.169.70|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:40 ERROR 404: Not Found.

