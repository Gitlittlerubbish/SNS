--2020-02-25 22:13:54--  https://www.promerica.com.sv/media/1229/reglamento.pdf%0D
Resolving www.promerica.com.sv (www.promerica.com.sv)... 45.60.154.167
Connecting to www.promerica.com.sv (www.promerica.com.sv)|45.60.154.167|:443... connected.
HTTP request sent, awaiting response... 403 Forbidden
2020-02-25 22:13:54 ERROR 403: Forbidden.

--2020-02-25 22:14:21--  https://www.promerica.com.sv/media/1229/reglamento.pdf%0D
Resolving www.promerica.com.sv (www.promerica.com.sv)... 45.60.154.167
Connecting to www.promerica.com.sv (www.promerica.com.sv)|45.60.154.167|:443... connected.
HTTP request sent, awaiting response... 403 Forbidden
2020-02-25 22:14:21 ERROR 403: Forbidden.

