--2020-02-25 22:13:55--  https://www.ugb.edu.sv/images/pdf/modeloeducativougb.pdf%0D
Resolving www.ugb.edu.sv (www.ugb.edu.sv)... 190.86.248.10
Connecting to www.ugb.edu.sv (www.ugb.edu.sv)|190.86.248.10|:443... connected.
HTTP request sent, awaiting response... 500 Internal Server Error
2020-02-25 22:13:56 ERROR 500: Internal Server Error.

--2020-02-25 22:14:21--  https://www.ugb.edu.sv/images/pdf/modeloeducativougb.pdf%0D
Resolving www.ugb.edu.sv (www.ugb.edu.sv)... 190.86.248.10
Connecting to www.ugb.edu.sv (www.ugb.edu.sv)|190.86.248.10|:443... connected.
HTTP request sent, awaiting response... 500 Internal Server Error
2020-02-25 22:14:23 ERROR 500: Internal Server Error.

