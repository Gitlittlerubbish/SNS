--2020-02-25 22:13:54--  http://santatecla.gob.sv/documentos/Servicios-Catastro.pdf%0D
Resolving santatecla.gob.sv (santatecla.gob.sv)... 192.254.190.129
Connecting to santatecla.gob.sv (santatecla.gob.sv)|192.254.190.129|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:55 ERROR 404: Not Found.

--2020-02-25 22:14:21--  http://santatecla.gob.sv/documentos/Servicios-Catastro.pdf%0D
Resolving santatecla.gob.sv (santatecla.gob.sv)... 192.254.190.129
Connecting to santatecla.gob.sv (santatecla.gob.sv)|192.254.190.129|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:21 ERROR 404: Not Found.

