--2020-03-02 03:23:56--  http://www.transparencia.gob.sv/institutions/isss/documents/7853/download
Resolving www.transparencia.gob.sv (www.transparencia.gob.sv)... 95.216.118.177
Connecting to www.transparencia.gob.sv (www.transparencia.gob.sv)|95.216.118.177|:80... connected.
HTTP request sent, awaiting response... 302 Found
Location: https://www.transparencia.gob.sv/institutions/isss/documents/7853/download [following]
--2020-03-02 03:23:57--  https://www.transparencia.gob.sv/institutions/isss/documents/7853/download
Connecting to www.transparencia.gob.sv (www.transparencia.gob.sv)|95.216.118.177|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 5.57M
    50K .......... .......... .......... .......... .......... 10.5M
   100K .......... .......... .......... .......... ..........  181M
   150K .......... .......... .......... .......... ..........  175M
   200K .......... .......... ........                         7.03M=0.2s

2020-03-02 03:23:57 (12.4 Mb/s) - ‘/dev/null’ saved [234015]

