--2020-03-02 03:23:57--  http://www.informacionpublicapgr.gob.sv/descargables/sia/normativa-internacional/Gestexto2.pdf
Resolving www.informacionpublicapgr.gob.sv (www.informacionpublicapgr.gob.sv)... 131.100.141.22
Connecting to www.informacionpublicapgr.gob.sv (www.informacionpublicapgr.gob.sv)|131.100.141.22|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 380590 (372K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 13%  993K 3s
    50K .......... .......... .......... .......... .......... 26% 2.85M 2s
   100K .......... .......... .......... .......... .......... 40% 50.9M 1s
   150K .......... .......... .......... .......... .......... 53% 3.07M 1s
   200K .......... .......... .......... .......... .......... 67% 50.1M 0s
   250K .......... .......... .......... .......... .......... 80%  108M 0s
   300K .......... .......... .......... .......... .......... 94% 3.12M 0s
   350K .......... .......... .                               100% 56.7M=0.8s

2020-03-02 03:23:58 (3.61 Mb/s) - ‘/dev/null’ saved [380590/380590]

