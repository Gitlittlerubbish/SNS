--2020-02-25 22:12:56--  https://prisma.org.sv/asset/documents/480%0D
Resolving prisma.org.sv (prisma.org.sv)... 192.241.239.186
Connecting to prisma.org.sv (prisma.org.sv)|192.241.239.186|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 1.38M
    50K .......... .......... .......... .......... .......... 2.78M
   100K .......... .......... .......... .......... ..........  999M
   150K .......... .......... .......... .......... .......... 2.79M
   200K .......... .......... .......... .......... ..........  781M
   250K .......... .......... .......... .......... ..........  859M
   300K .......... .......... .                                2.33G=0.6s

2020-02-25 22:12:58 (4.45 Mb/s) - ‘/dev/null’ saved [329595]

--2020-02-25 22:12:58--  https://prisma.org.sv/asset/documents/480%0D
Resolving prisma.org.sv (prisma.org.sv)... 192.241.239.186
Connecting to prisma.org.sv (prisma.org.sv)|192.241.239.186|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 1.40M
    50K .......... .......... .......... .......... .......... 2.82M
   100K .......... .......... .......... .......... ..........  606M
   150K .......... .......... .......... .......... .......... 2.82M
   200K .......... .......... .......... .......... .......... 1.02G
   250K .......... .......... .......... .......... .......... 1.28G
   300K .......... .......... .                                1.61G=0.6s

2020-02-25 22:12:59 (4.52 Mb/s) - ‘/dev/null’ saved [329595]

--2020-02-25 22:13:32--  https://prisma.org.sv/asset/documents/480%0D
Resolving prisma.org.sv (prisma.org.sv)... 192.241.239.186
Connecting to prisma.org.sv (prisma.org.sv)|192.241.239.186|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 1.42M
    50K .......... .......... .......... .......... .......... 2.83M
   100K .......... .......... .......... .......... ..........  353M
   150K .......... .......... .......... .......... .......... 2.86M
   200K .......... .......... .......... .......... .......... 1.22G
   250K .......... .......... .......... .......... ..........  981M
   300K .......... .......... .                                 878M=0.6s

2020-02-25 22:13:33 (4.56 Mb/s) - ‘/dev/null’ saved [329595]

--2020-02-25 22:13:33--  https://prisma.org.sv/asset/documents/480%0D
Resolving prisma.org.sv (prisma.org.sv)... 192.241.239.186
Connecting to prisma.org.sv (prisma.org.sv)|192.241.239.186|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 1.43M
    50K .......... .......... .......... .......... .......... 2.86M
   100K .......... .......... .......... .......... ..........  610M
   150K .......... .......... .......... .......... .......... 2.86M
   200K .......... .......... .......... .......... .......... 1.20G
   250K .......... .......... .......... .......... .......... 1.59G
   300K .......... .......... .                                1.47G=0.6s

2020-02-25 22:13:34 (4.59 Mb/s) - ‘/dev/null’ saved [329595]

