--2020-02-25 22:12:47--  https://www.mined.gob.sv/sexualidad/Media.pdf%0D
Resolving www.mined.gob.sv (www.mined.gob.sv)... 168.243.116.34
Connecting to www.mined.gob.sv (www.mined.gob.sv)|168.243.116.34|:443... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:12:47 ERROR 404: Not Found.

--2020-02-25 22:13:25--  https://www.mined.gob.sv/sexualidad/Media.pdf%0D
Resolving www.mined.gob.sv (www.mined.gob.sv)... 168.243.116.34
Connecting to www.mined.gob.sv (www.mined.gob.sv)|168.243.116.34|:443... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:25 ERROR 404: Not Found.

