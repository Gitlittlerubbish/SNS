--2020-02-25 22:12:43--  http://www.yamaha-motor.com.sv/home/storage/documents/QvbsNSQyqeaYdfIBTUK5KxEZCJEDABeZlmzDjQXM.pdf%0D
Resolving www.yamaha-motor.com.sv (www.yamaha-motor.com.sv)... 72.47.228.69
Connecting to www.yamaha-motor.com.sv (www.yamaha-motor.com.sv)|72.47.228.69|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:12:45 ERROR 404: Not Found.

--2020-02-25 22:13:23--  http://www.yamaha-motor.com.sv/home/storage/documents/QvbsNSQyqeaYdfIBTUK5KxEZCJEDABeZlmzDjQXM.pdf%0D
Resolving www.yamaha-motor.com.sv (www.yamaha-motor.com.sv)... 72.47.228.69
Connecting to www.yamaha-motor.com.sv (www.yamaha-motor.com.sv)|72.47.228.69|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:24 ERROR 404: Not Found.

