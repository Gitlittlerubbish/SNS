--2020-02-25 22:13:34--  http://www.grupoacc.com.sv/Files/DEC_160.pdf%0D
Resolving www.grupoacc.com.sv (www.grupoacc.com.sv)... 192.185.148.210
Connecting to www.grupoacc.com.sv (www.grupoacc.com.sv)|192.185.148.210|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:35 ERROR 404: Not Found.

--2020-02-25 22:14:08--  http://www.grupoacc.com.sv/Files/DEC_160.pdf%0D
Resolving www.grupoacc.com.sv (www.grupoacc.com.sv)... 192.185.148.210
Connecting to www.grupoacc.com.sv (www.grupoacc.com.sv)|192.185.148.210|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:08 ERROR 404: Not Found.

