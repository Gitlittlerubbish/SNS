--2020-02-25 22:12:51--  http://www.islam.org.sv/biblioteca/El_Verdadero_Mensaje_de_Jesucristo.pdf%0D
Resolving www.islam.org.sv (www.islam.org.sv)... failed: Name or service not known.
wget: unable to resolve host address ‘www.islam.org.sv’
--2020-02-25 22:13:28--  http://www.islam.org.sv/biblioteca/El_Verdadero_Mensaje_de_Jesucristo.pdf%0D
Resolving www.islam.org.sv (www.islam.org.sv)... failed: Name or service not known.
wget: unable to resolve host address ‘www.islam.org.sv’
