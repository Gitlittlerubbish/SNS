--2020-03-02 03:24:27--  http://www.snet.gob.sv/Geologia/DeslavePicacho.pdf
Resolving www.snet.gob.sv (www.snet.gob.sv)... 190.5.148.229, 170.0.177.4
Connecting to www.snet.gob.sv (www.snet.gob.sv)|190.5.148.229|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 740013 (723K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  6% 1.46M 4s
    50K .......... .......... .......... .......... .......... 13% 3.02M 3s
   100K .......... .......... .......... .......... .......... 20% 55.6M 2s
   150K .......... .......... .......... .......... .......... 27% 81.2M 1s
   200K .......... .......... .......... .......... .......... 34% 3.03M 1s
   250K .......... .......... .......... .......... .......... 41% 45.3M 1s
   300K .......... .......... .......... .......... .......... 48% 3.31M 1s
   350K .......... .......... .......... .......... .......... 55% 49.4M 1s
   400K .......... .......... .......... .......... .......... 62% 2.63M 1s
   450K .......... .......... .......... .......... .......... 69% 21.6M 0s
   500K .......... .......... .......... .......... .......... 76% 1.39G 0s
   550K .......... .......... .......... .......... .......... 83% 1.46G 0s
   600K .......... .......... .......... .......... .......... 89% 1.31G 0s
   650K .......... .......... .......... .......... .......... 96% 3.49M 0s
   700K .......... .......... ..                              100% 10.4M=1.0s

2020-03-02 03:24:28 (5.83 Mb/s) - ‘/dev/null’ saved [740013/740013]

