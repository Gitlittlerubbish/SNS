--2020-03-02 03:24:31--  http://prisma.org.sv/asset/documents/480
Resolving prisma.org.sv (prisma.org.sv)... 192.241.239.186
Connecting to prisma.org.sv (prisma.org.sv)|192.241.239.186|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: https://prisma.org.sv/asset/documents/480 [following]
--2020-03-02 03:24:31--  https://prisma.org.sv/asset/documents/480
Connecting to prisma.org.sv (prisma.org.sv)|192.241.239.186|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 1.36M
    50K .......... .......... .......... .......... .......... 2.77M
   100K .......... .......... .......... .......... ..........  103M
   150K .......... .......... .......... .......... .......... 2.84M
   200K .......... .......... .......... .......... ..........  119M
   250K .......... .......... .......... .......... .......... 80.1M
   300K .......... .......... .                                40.4M=0.6s

2020-03-02 03:24:32 (4.32 Mb/s) - ‘/dev/null’ saved [329595]

