--2020-02-25 22:14:04--  https://defensoria.gob.sv/wp-content/uploads/2015/04/92-DO_NSO_67_32_03_03control_visual.pdf%0D
Resolving defensoria.gob.sv (defensoria.gob.sv)... 190.5.140.226
Connecting to defensoria.gob.sv (defensoria.gob.sv)|190.5.140.226|:443... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: https://www.defensoria.gob.sv/wp-content/uploads/2015/04/92-DO_NSO_67_32_03_03control_visual.pdf [following]
--2020-02-25 22:14:07--  https://www.defensoria.gob.sv/wp-content/uploads/2015/04/92-DO_NSO_67_32_03_03control_visual.pdf
Resolving www.defensoria.gob.sv (www.defensoria.gob.sv)... 190.5.140.226
Connecting to www.defensoria.gob.sv (www.defensoria.gob.sv)|190.5.140.226|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: 1076990 (1.0M) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  4% 1.48M 6s
    50K .......... .......... .......... .......... ..........  9% 1.59M 5s
   100K .......... .......... .......... .......... .......... 14% 97.8M 3s
   150K .......... .......... .......... .......... .......... 19% 3.10M 3s
   200K .......... .......... .......... .......... .......... 23% 95.7M 2s
   250K .......... .......... .......... .......... .......... 28% 3.16M 2s
   300K .......... .......... .......... .......... .......... 33% 97.6M 2s
   350K .......... .......... .......... .......... .......... 38% 95.0M 1s
   400K .......... .......... .......... .......... .......... 42% 3.25M 1s
   450K .......... .......... .......... .......... .......... 47% 95.3M 1s
   500K .......... .......... .......... .......... .......... 52% 95.1M 1s
   550K .......... .......... .......... .......... .......... 57% 84.9M 1s
   600K .......... .......... .......... .......... .......... 61% 89.4M 1s
   650K .......... .......... .......... .......... .......... 66% 3.51M 1s
   700K .......... .......... .......... .......... .......... 71% 89.8M 0s
   750K .......... .......... .......... .......... .......... 76% 94.2M 0s
   800K .......... .......... .......... .......... .......... 80% 71.6M 0s
   850K .......... .......... .......... .......... .......... 85% 94.6M 0s
   900K .......... .......... .......... .......... .......... 90% 94.1M 0s
   950K .......... .......... .......... .......... .......... 95% 3.83M 0s
  1000K .......... .......... .......... .......... .......... 99%  112M 0s
  1050K .                                                     100% 28640G=1.2s

2020-02-25 22:14:09 (7.13 Mb/s) - ‘/dev/null’ saved [1076990/1076990]

--2020-02-25 22:14:09--  https://defensoria.gob.sv/wp-content/uploads/2015/04/92-DO_NSO_67_32_03_03control_visual.pdf%0D
Resolving defensoria.gob.sv (defensoria.gob.sv)... 190.5.140.226
Connecting to defensoria.gob.sv (defensoria.gob.sv)|190.5.140.226|:443... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: https://www.defensoria.gob.sv/wp-content/uploads/2015/04/92-DO_NSO_67_32_03_03control_visual.pdf [following]
--2020-02-25 22:14:12--  https://www.defensoria.gob.sv/wp-content/uploads/2015/04/92-DO_NSO_67_32_03_03control_visual.pdf
Resolving www.defensoria.gob.sv (www.defensoria.gob.sv)... 190.5.140.226
Connecting to www.defensoria.gob.sv (www.defensoria.gob.sv)|190.5.140.226|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: 1076990 (1.0M) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  4% 1.05M 8s
    50K .......... .......... .......... .......... ..........  9% 3.13M 5s
   100K .......... .......... .......... .......... .......... 14% 3.18M 4s
   150K .......... .......... .......... .......... .......... 19% 90.7M 3s
   200K .......... .......... .......... .......... .......... 23% 3.25M 3s
   250K .......... .......... .......... .......... .......... 28% 97.4M 2s
   300K .......... .......... .......... .......... .......... 33% 94.6M 2s
   350K .......... .......... .......... .......... .......... 38% 3.35M 1s
   400K .......... .......... .......... .......... .......... 42% 72.5M 1s
   450K .......... .......... .......... .......... .......... 47% 94.1M 1s
   500K .......... .......... .......... .......... .......... 52% 92.8M 1s
   550K .......... .......... .......... .......... .......... 57% 3.53M 1s
   600K .......... .......... .......... .......... .......... 61% 95.9M 1s
   650K .......... .......... .......... .......... .......... 66% 89.7M 1s
   700K .......... .......... .......... .......... .......... 71% 95.3M 0s
   750K .......... .......... .......... .......... .......... 76% 93.0M 0s
   800K .......... .......... .......... .......... .......... 80% 67.0M 0s
   850K .......... .......... .......... .......... .......... 85% 3.85M 0s
   900K .......... .......... .......... .......... .......... 90% 98.1M 0s
   950K .......... .......... .......... .......... .......... 95% 88.0M 0s
  1000K .......... .......... .......... .......... .......... 99%  105M 0s
  1050K .                                                     100% 28640G=1.2s

2020-02-25 22:14:13 (7.27 Mb/s) - ‘/dev/null’ saved [1076990/1076990]

--2020-02-25 22:14:30--  https://defensoria.gob.sv/wp-content/uploads/2015/04/92-DO_NSO_67_32_03_03control_visual.pdf%0D
Resolving defensoria.gob.sv (defensoria.gob.sv)... 190.5.140.226
Connecting to defensoria.gob.sv (defensoria.gob.sv)|190.5.140.226|:443... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: https://www.defensoria.gob.sv/wp-content/uploads/2015/04/92-DO_NSO_67_32_03_03control_visual.pdf [following]
--2020-02-25 22:14:32--  https://www.defensoria.gob.sv/wp-content/uploads/2015/04/92-DO_NSO_67_32_03_03control_visual.pdf
Resolving www.defensoria.gob.sv (www.defensoria.gob.sv)... 190.5.140.226
Connecting to www.defensoria.gob.sv (www.defensoria.gob.sv)|190.5.140.226|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: 1076990 (1.0M) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  4% 1.36M 6s
    50K .......... .......... .......... .......... ..........  9% 4.40M 4s
   100K .......... .......... .......... .......... .......... 14% 3.18M 3s
   150K .......... .......... .......... .......... .......... 19% 90.2M 2s
   200K .......... .......... .......... .......... .......... 23% 3.27M 2s
   250K .......... .......... .......... .......... .......... 28% 96.9M 2s
   300K .......... .......... .......... .......... .......... 33% 95.5M 1s
   350K .......... .......... .......... .......... .......... 38% 6.02M 1s
   400K .......... .......... .......... .......... .......... 42% 7.27M 1s
   450K .......... .......... .......... .......... .......... 47% 84.1M 1s
   500K .......... .......... .......... .......... .......... 52% 96.2M 1s
   550K .......... .......... .......... .......... .......... 57% 80.5M 1s
   600K .......... .......... .......... .......... .......... 61% 96.6M 0s
   650K .......... .......... .......... .......... .......... 66% 21.8M 0s
   700K .......... .......... .......... .......... .......... 71% 4.53M 0s
   750K .......... .......... .......... .......... .......... 76% 95.2M 0s
   800K .......... .......... .......... .......... .......... 80% 65.8M 0s
   850K .......... .......... .......... .......... .......... 85% 83.2M 0s
   900K .......... .......... .......... .......... .......... 90% 86.5M 0s
   950K .......... .......... .......... .......... .......... 95% 95.5M 0s
  1000K .......... .......... .......... .......... .......... 99%  105M 0s
  1050K .                                                     100% 28640G=0.9s

2020-02-25 22:14:34 (9.16 Mb/s) - ‘/dev/null’ saved [1076990/1076990]

--2020-02-25 22:14:34--  https://defensoria.gob.sv/wp-content/uploads/2015/04/92-DO_NSO_67_32_03_03control_visual.pdf%0D
Resolving defensoria.gob.sv (defensoria.gob.sv)... 190.5.140.226
Connecting to defensoria.gob.sv (defensoria.gob.sv)|190.5.140.226|:443... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: https://www.defensoria.gob.sv/wp-content/uploads/2015/04/92-DO_NSO_67_32_03_03control_visual.pdf [following]
--2020-02-25 22:14:36--  https://www.defensoria.gob.sv/wp-content/uploads/2015/04/92-DO_NSO_67_32_03_03control_visual.pdf
Resolving www.defensoria.gob.sv (www.defensoria.gob.sv)... 190.5.140.226
Connecting to www.defensoria.gob.sv (www.defensoria.gob.sv)|190.5.140.226|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: 1076990 (1.0M) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  4% 1.06M 8s
    50K .......... .......... .......... .......... ..........  9% 3.18M 5s
   100K .......... .......... .......... .......... .......... 14% 89.6M 3s
   150K .......... .......... .......... .......... .......... 19% 3.22M 3s
   200K .......... .......... .......... .......... .......... 23% 90.3M 2s
   250K .......... .......... .......... .......... .......... 28% 3.31M 2s
   300K .......... .......... .......... .......... .......... 33% 94.2M 2s
   350K .......... .......... .......... .......... .......... 38% 88.7M 1s
   400K .......... .......... .......... .......... .......... 42% 3.39M 1s
   450K .......... .......... .......... .......... .......... 47% 86.9M 1s
   500K .......... .......... .......... .......... .......... 52% 84.6M 1s
   550K .......... .......... .......... .......... .......... 57% 89.4M 1s
   600K .......... .......... .......... .......... .......... 61% 3.65M 1s
   650K .......... .......... .......... .......... .......... 66% 94.7M 1s
   700K .......... .......... .......... .......... .......... 71% 87.3M 0s
   750K .......... .......... .......... .......... .......... 76% 94.8M 0s
   800K .......... .......... .......... .......... .......... 80% 71.3M 0s
   850K .......... .......... .......... .......... .......... 85% 84.5M 0s
   900K .......... .......... .......... .......... .......... 90% 3.98M 0s
   950K .......... .......... .......... .......... .......... 95% 94.0M 0s
  1000K .......... .......... .......... .......... .......... 99%  106M 0s
  1050K .                                                     100% 28640G=1.2s

2020-02-25 22:14:38 (7.39 Mb/s) - ‘/dev/null’ saved [1076990/1076990]

