--2020-02-25 22:12:53--  http://www.sc.gob.sv/uploads/est_24_inf.pdf%0D
Resolving www.sc.gob.sv (www.sc.gob.sv)... 190.5.133.234
Connecting to www.sc.gob.sv (www.sc.gob.sv)|190.5.133.234|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:12:54 ERROR 404: Not Found.

--2020-02-25 22:13:29--  http://www.sc.gob.sv/uploads/est_24_inf.pdf%0D
Resolving www.sc.gob.sv (www.sc.gob.sv)... 190.5.133.234
Connecting to www.sc.gob.sv (www.sc.gob.sv)|190.5.133.234|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:30 ERROR 404: Not Found.

