--2020-03-02 03:26:05--  http://www.salud.gob.sv/archivos/vigi_epide2019/Calendario_Epidemiologico_2019.pdf
Resolving www.salud.gob.sv (www.salud.gob.sv)... 190.86.223.123
Connecting to www.salud.gob.sv (www.salud.gob.sv)|190.86.223.123|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 153378 (150K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 33% 1.57M 1s
    50K .......... .......... .......... .......... .......... 66% 3.01M 0s
   100K .......... .......... .......... .......... ......... 100% 1.35G=0.4s

2020-03-02 03:26:06 (3.09 Mb/s) - ‘/dev/null’ saved [153378/153378]

