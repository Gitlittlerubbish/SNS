--2020-03-02 03:25:35--  http://www.mh.gob.sv/downloads/pdf/PMHDC8306.pdf
Resolving www.mh.gob.sv (www.mh.gob.sv)... 190.5.131.13, 190.57.24.24
Connecting to www.mh.gob.sv (www.mh.gob.sv)|190.5.131.13|:80... connected.
HTTP request sent, awaiting response... 302 Moved Temporarily
Location: https://www.mh.gob.sv/downloads/pdf/PMHDC8306.pdf [following]
--2020-03-02 03:25:36--  https://www.mh.gob.sv/downloads/pdf/PMHDC8306.pdf
Connecting to www.mh.gob.sv (www.mh.gob.sv)|190.5.131.13|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: 553570 (541K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  9% 1.46M 3s
    50K .......... .......... .......... .......... .......... 18% 2.75M 2s
   100K .......... .......... .......... .......... .......... 27% 2.81M 1s
   150K .......... .......... .......... .......... .......... 36% 2.84M 1s
   200K .......... .......... .......... .......... .......... 46% 1.76M 1s
   250K .......... .......... .......... .......... .......... 55% 2.18M 1s
   300K .......... .......... .......... .......... .......... 64% 2.77M 1s
   350K .......... .......... .......... .......... .......... 73% 2.90M 1s
   400K .......... .......... .......... .......... .......... 83% 1.73M 0s
   450K .......... .......... .......... .......... .......... 92% 2.17M 0s
   500K .......... .......... .......... ..........           100% 2.35M=2.0s

2020-03-02 03:25:38 (2.22 Mb/s) - ‘/dev/null’ saved [553570/553570]

