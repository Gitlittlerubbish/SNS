--2020-03-02 03:25:04--  http://thyssenkrupp.com.sv/noticia/download/763/
Resolving thyssenkrupp.com.sv (thyssenkrupp.com.sv)... 186.202.143.17
Connecting to thyssenkrupp.com.sv (thyssenkrupp.com.sv)|186.202.143.17|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: https://thyssenkrupp.com.sv/noticia/download/763/ [following]
--2020-03-02 03:25:05--  https://thyssenkrupp.com.sv/noticia/download/763/
Connecting to thyssenkrupp.com.sv (thyssenkrupp.com.sv)|186.202.143.17|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: 1282642 (1.2M) [application/download]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  3%  778K 13s
    50K .......... .......... .......... .......... ..........  7% 1.56M 9s
   100K .......... .......... .......... .......... .......... 11%  123M 6s
   150K .......... .......... .......... .......... .......... 15% 1.56M 6s
   200K .......... .......... .......... .......... .......... 19% 1.56M 5s
   250K .......... .......... .......... .......... .......... 23% 1.56M 5s
   300K .......... .......... .......... .......... .......... 27% 1.58M 5s
   350K .......... .......... .......... .......... .......... 31% 60.3M 4s
   400K .......... .......... .......... .......... .......... 35% 1.56M 4s
   450K .......... .......... .......... .......... .......... 39% 1.56M 4s
   500K .......... .......... .......... .......... .......... 43% 1.55M 3s
   550K .......... .......... .......... .......... .......... 47% 4.20M 3s
   600K .......... .......... .......... .......... .......... 51% 2.47M 3s
   650K .......... .......... .......... .......... .......... 55% 1.56M 2s
   700K .......... .......... .......... .......... .......... 59% 1.56M 2s
   750K .......... .......... .......... .......... .......... 63% 1.55M 2s
   800K .......... .......... .......... .......... .......... 67% 1.62M 2s
   850K .......... .......... .......... .......... .......... 71% 3.74M 2s
   900K .......... .......... .......... .......... .......... 75% 2.47M 1s
   950K .......... .......... .......... .......... .......... 79% 1.56M 1s
  1000K .......... .......... .......... .......... .......... 83% 1.63M 1s
  1050K .......... .......... .......... .......... .......... 87% 1.98M 1s
  1100K .......... .......... .......... .......... .......... 91% 5.79M 0s
  1150K .......... .......... .......... .......... .......... 95% 1.58M 0s
  1200K .......... .......... .......... .......... .......... 99% 1.56M 0s
  1250K ..                                                    100%  181M=5.5s

2020-03-02 03:25:12 (1.86 Mb/s) - ‘/dev/null’ saved [1282642/1282642]

