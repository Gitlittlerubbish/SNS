--2020-03-02 03:26:17--  http://ui.usonsonate.edu.sv/papers/DIRECTORES_EXITOSOS.pdf
Resolving ui.usonsonate.edu.sv (ui.usonsonate.edu.sv)... 66.113.161.172
Connecting to ui.usonsonate.edu.sv (ui.usonsonate.edu.sv)|66.113.161.172|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 1707851 (1.6M) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  2% 1.76M 8s
    50K .......... .......... .......... .......... ..........  5% 3.53M 5s
   100K .......... .......... .......... .......... ..........  8% 3.43M 5s
   150K .......... .......... .......... .......... .......... 11% 3.59M 4s
   200K .......... .......... .......... .......... .......... 14% 90.7M 3s
   250K .......... .......... .......... .......... .......... 17% 3.70M 3s
   300K .......... .......... .......... .......... .......... 20% 99.7M 3s
   350K .......... .......... .......... .......... .......... 23%  107M 2s
   400K .......... .......... .......... .......... .......... 26% 3.79M 2s
   450K .......... .......... .......... .......... .......... 29% 55.0M 2s
   500K .......... .......... .......... .......... .......... 32%  138M 2s
   550K .......... .......... .......... .......... .......... 35%  154M 1s
   600K .......... .......... .......... .......... .......... 38% 70.1M 1s
   650K .......... .......... .......... .......... .......... 41% 4.06M 1s
   700K .......... .......... .......... .......... .......... 44% 83.6M 1s
   750K .......... .......... .......... .......... .......... 47% 97.6M 1s
   800K .......... .......... .......... .......... .......... 50% 82.9M 1s
   850K .......... .......... .......... .......... .......... 53%  128M 1s
   900K .......... .......... .......... .......... .......... 56% 4.16M 1s
   950K .......... .......... .......... .......... .......... 59% 72.3M 1s
  1000K .......... .......... .......... .......... .......... 62%  173M 1s
  1050K .......... .......... .......... .......... .......... 65%  116M 1s
  1100K .......... .......... .......... .......... .......... 68% 56.9M 0s
  1150K .......... .......... .......... .......... .......... 71%  135M 0s
  1200K .......... .......... .......... .......... .......... 74%  197M 0s
  1250K .......... .......... .......... .......... .......... 77% 53.1M 0s
  1300K .......... .......... .......... .......... .......... 80% 4.71M 0s
  1350K .......... .......... .......... .......... .......... 83% 96.4M 0s
  1400K .......... .......... .......... .......... .......... 86% 52.6M 0s
  1450K .......... .......... .......... .......... .......... 89% 53.7M 0s
  1500K .......... .......... .......... .......... .......... 92%  168M 0s
  1550K .......... .......... .......... .......... .......... 95% 56.0M 0s
  1600K .......... .......... .......... .......... .......... 98%  301M 0s
  1650K .......... .......                                    100% 46.9M=1.2s

2020-03-02 03:26:19 (11.4 Mb/s) - ‘/dev/null’ saved [1707851/1707851]

