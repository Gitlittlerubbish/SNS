--2020-02-25 22:12:43--  http://www.informacionpublicapgr.gob.sv/descargables/sia/normativa-internacional/Gestexto2.pdf%0D
Resolving www.informacionpublicapgr.gob.sv (www.informacionpublicapgr.gob.sv)... 131.100.141.22
Connecting to www.informacionpublicapgr.gob.sv (www.informacionpublicapgr.gob.sv)|131.100.141.22|:80... connected.
HTTP request sent, awaiting response... 403 Forbidden
2020-02-25 22:12:43 ERROR 403: Forbidden.

--2020-02-25 22:13:23--  http://www.informacionpublicapgr.gob.sv/descargables/sia/normativa-internacional/Gestexto2.pdf%0D
Resolving www.informacionpublicapgr.gob.sv (www.informacionpublicapgr.gob.sv)... 131.100.141.22
Connecting to www.informacionpublicapgr.gob.sv (www.informacionpublicapgr.gob.sv)|131.100.141.22|:80... connected.
HTTP request sent, awaiting response... 403 Forbidden
2020-02-25 22:13:23 ERROR 403: Forbidden.

