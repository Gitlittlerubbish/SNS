--2020-03-02 03:24:20--  http://www.sc.gob.sv/uploads/est_24_inf.pdf
Resolving www.sc.gob.sv (www.sc.gob.sv)... 190.5.133.234
Connecting to www.sc.gob.sv (www.sc.gob.sv)|190.5.133.234|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 5150630 (4.9M) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  0% 1.49M 27s
    50K .......... .......... .......... .......... ..........  1% 3.15M 20s
   100K .......... .......... .......... .......... ..........  2% 8.30M 15s
   150K .......... .......... .......... .......... ..........  3% 8.84M 12s
   200K .......... .......... .......... .......... ..........  4% 5.52M 11s
   250K .......... .......... .......... .......... ..........  5% 8.20M 10s
   300K .......... .......... .......... .......... ..........  6% 7.13M 9s
   350K .......... .......... .......... .......... ..........  7% 8.03M 8s
   400K .......... .......... .......... .......... ..........  8% 8.18M 8s
   450K .......... .......... .......... .......... ..........  9% 8.30M 8s
   500K .......... .......... .......... .......... .......... 10% 8.00M 7s
   550K .......... .......... .......... .......... .......... 11% 8.23M 7s
   600K .......... .......... .......... .......... .......... 12% 8.20M 7s
   650K .......... .......... .......... .......... .......... 13% 8.21M 6s
   700K .......... .......... .......... .......... .......... 14% 8.05M 6s
   750K .......... .......... .......... .......... .......... 15% 8.05M 6s
   800K .......... .......... .......... .......... .......... 16% 8.69M 6s
   850K .......... .......... .......... .......... .......... 17% 8.09M 6s
   900K .......... .......... .......... .......... .......... 18% 7.77M 6s
   950K .......... .......... .......... .......... .......... 19% 8.33M 5s
  1000K .......... .......... .......... .......... .......... 20% 8.13M 5s
  1050K .......... .......... .......... .......... .......... 21% 7.95M 5s
  1100K .......... .......... .......... .......... .......... 22% 8.48M 5s
  1150K .......... .......... .......... .......... .......... 23% 8.24M 5s
  1200K .......... .......... .......... .......... .......... 24% 8.34M 5s
  1250K .......... .......... .......... .......... .......... 25% 7.81M 5s
  1300K .......... .......... .......... .......... .......... 26% 8.52M 5s
  1350K .......... .......... .......... .......... .......... 27% 8.15M 4s
  1400K .......... .......... .......... .......... .......... 28% 7.99M 4s
  1450K .......... .......... .......... .......... .......... 29% 8.35M 4s
  1500K .......... .......... .......... .......... .......... 30% 4.06M 4s
  1550K .......... .......... .......... .......... .......... 31%  154M 4s
  1600K .......... .......... .......... .......... .......... 32% 8.50M 4s
  1650K .......... .......... .......... .......... .......... 33% 8.19M 4s
  1700K .......... .......... .......... .......... .......... 34% 8.26M 4s
  1750K .......... .......... .......... .......... .......... 35% 7.97M 4s
  1800K .......... .......... .......... .......... .......... 36% 8.40M 4s
  1850K .......... .......... .......... .......... .......... 37% 8.16M 4s
  1900K .......... .......... .......... .......... .......... 38% 8.48M 4s
  1950K .......... .......... .......... .......... .......... 39% 8.23M 4s
  2000K .......... .......... .......... .......... .......... 40% 7.84M 3s
  2050K .......... .......... .......... .......... .......... 41% 8.02M 3s
  2100K .......... .......... .......... .......... .......... 42% 8.38M 3s
  2150K .......... .......... .......... .......... .......... 43% 8.28M 3s
  2200K .......... .......... .......... .......... .......... 44% 8.00M 3s
  2250K .......... .......... .......... .......... .......... 45% 8.30M 3s
  2300K .......... .......... .......... .......... .......... 46% 8.16M 3s
  2350K .......... .......... .......... .......... .......... 47% 7.93M 3s
  2400K .......... .......... .......... .......... .......... 48% 8.11M 3s
  2450K .......... .......... .......... .......... .......... 49% 8.24M 3s
  2500K .......... .......... .......... .......... .......... 50% 8.56M 3s
  2550K .......... .......... .......... .......... .......... 51% 8.12M 3s
  2600K .......... .......... .......... .......... .......... 52% 8.29M 3s
  2650K .......... .......... .......... .......... .......... 53% 7.96M 3s
  2700K .......... .......... .......... .......... .......... 54% 8.49M 3s
  2750K .......... .......... .......... .......... .......... 55% 8.23M 2s
  2800K .......... .......... .......... .......... .......... 56% 8.06M 2s
  2850K .......... .......... .......... .......... .......... 57% 7.81M 2s
  2900K .......... .......... .......... .......... .......... 58% 8.48M 2s
  2950K .......... .......... .......... .......... .......... 59% 8.08M 2s
  3000K .......... .......... .......... .......... .......... 60% 7.97M 2s
  3050K .......... .......... .......... .......... .......... 61% 8.32M 2s
  3100K .......... .......... .......... .......... .......... 62% 8.20M 2s
  3150K .......... .......... .......... .......... .......... 63% 8.49M 2s
  3200K .......... .......... .......... .......... .......... 64% 8.13M 2s
  3250K .......... .......... .......... .......... .......... 65% 8.02M 2s
  3300K .......... .......... .......... .......... .......... 66% 7.94M 2s
  3350K .......... .......... .......... .......... .......... 67% 8.23M 2s
  3400K .......... .......... .......... .......... .......... 68% 8.44M 2s
  3450K .......... .......... .......... .......... .......... 69% 8.27M 2s
  3500K .......... .......... .......... .......... .......... 70% 8.36M 2s
  3550K .......... .......... .......... .......... .......... 71% 8.06M 2s
  3600K .......... .......... .......... .......... .......... 72% 7.78M 2s
  3650K .......... .......... .......... .......... .......... 73% 8.34M 1s
  3700K .......... .......... .......... .......... .......... 74% 8.20M 1s
  3750K .......... .......... .......... .......... .......... 75% 8.06M 1s
  3800K .......... .......... .......... .......... .......... 76% 8.25M 1s
  3850K .......... .......... .......... .......... .......... 77% 8.54M 1s
  3900K .......... .......... .......... .......... .......... 78% 7.55M 1s
  3950K .......... .......... .......... .......... .......... 79% 8.51M 1s
  4000K .......... .......... .......... .......... .......... 80% 7.95M 1s
  4050K .......... .......... .......... .......... .......... 81% 8.65M 1s
  4100K .......... .......... .......... .......... .......... 82% 7.80M 1s
  4150K .......... .......... .......... .......... .......... 83% 8.19M 1s
  4200K .......... .......... .......... .......... .......... 84% 8.38M 1s
  4250K .......... .......... .......... .......... .......... 85% 8.05M 1s
  4300K .......... .......... .......... .......... .......... 86% 8.46M 1s
  4350K .......... .......... .......... .......... .......... 87% 8.43M 1s
  4400K .......... .......... .......... .......... .......... 88% 8.00M 1s
  4450K .......... .......... .......... .......... .......... 89% 7.94M 1s
  4500K .......... .......... .......... .......... .......... 90% 8.19M 1s
  4550K .......... .......... .......... .......... .......... 91% 8.00M 0s
  4600K .......... .......... .......... .......... .......... 92% 8.26M 0s
  4650K .......... .......... .......... .......... .......... 93% 8.35M 0s
  4700K .......... .......... .......... .......... .......... 94% 7.96M 0s
  4750K .......... .......... .......... .......... .......... 95% 8.59M 0s
  4800K .......... .......... .......... .......... .......... 96% 7.95M 0s
  4850K .......... .......... .......... .......... .......... 97% 8.70M 0s
  4900K .......... .......... .......... .......... .......... 98% 7.92M 0s
  4950K .......... .......... .......... .......... .......... 99% 8.03M 0s
  5000K .......... .......... .........                       100% 7.88M=5.4s

2020-03-02 03:24:26 (7.67 Mb/s) - ‘/dev/null’ saved [5150630/5150630]

