--2020-02-25 22:12:37--  http://www.uca.edu.sv/-pDIq89%0D
Resolving www.uca.edu.sv (www.uca.edu.sv)... 201.131.110.4
Connecting to www.uca.edu.sv (www.uca.edu.sv)|201.131.110.4|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 290 [text/html]
Saving to: ‘/dev/null’

     0K                                                       100%  670M=0s

2020-02-25 22:12:40 (670 Mb/s) - ‘/dev/null’ saved [290/290]

--2020-02-25 22:12:40--  http://www.uca.edu.sv/-pDIq89%0D
Resolving www.uca.edu.sv (www.uca.edu.sv)... 201.131.110.4
Connecting to www.uca.edu.sv (www.uca.edu.sv)|201.131.110.4|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 290 [text/html]
Saving to: ‘/dev/null’

     0K                                                       100%  315M=0s

2020-02-25 22:12:41 (315 Mb/s) - ‘/dev/null’ saved [290/290]

--2020-02-25 22:12:41--  http://www.uca.edu.sv/-1DUgTd%0D
Resolving www.uca.edu.sv (www.uca.edu.sv)... 201.131.110.4
Connecting to www.uca.edu.sv (www.uca.edu.sv)|201.131.110.4|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 274 [text/html]
Saving to: ‘/dev/null’

     0K                                                       100%  595M=0s

2020-02-25 22:12:41 (595 Mb/s) - ‘/dev/null’ saved [274/274]

--2020-02-25 22:12:41--  http://www.uca.edu.sv/-1DUgTd%0D
Resolving www.uca.edu.sv (www.uca.edu.sv)... 201.131.110.4
Connecting to www.uca.edu.sv (www.uca.edu.sv)|201.131.110.4|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 274 [text/html]
Saving to: ‘/dev/null’

     0K                                                       100%  585M=0s

2020-02-25 22:12:41 (585 Mb/s) - ‘/dev/null’ saved [274/274]

--2020-02-25 22:13:21--  http://www.uca.edu.sv/-pDIq89%0D
Resolving www.uca.edu.sv (www.uca.edu.sv)... 201.131.110.4
Connecting to www.uca.edu.sv (www.uca.edu.sv)|201.131.110.4|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 290 [text/html]
Saving to: ‘/dev/null’

     0K                                                       100%  311M=0s

2020-02-25 22:13:21 (311 Mb/s) - ‘/dev/null’ saved [290/290]

--2020-02-25 22:13:21--  http://www.uca.edu.sv/-pDIq89%0D
Resolving www.uca.edu.sv (www.uca.edu.sv)... 201.131.110.4
Connecting to www.uca.edu.sv (www.uca.edu.sv)|201.131.110.4|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 290 [text/html]
Saving to: ‘/dev/null’

     0K                                                       100%  112M=0s

2020-02-25 22:13:22 (112 Mb/s) - ‘/dev/null’ saved [290/290]

--2020-02-25 22:13:22--  http://www.uca.edu.sv/-1DUgTd%0D
Resolving www.uca.edu.sv (www.uca.edu.sv)... 201.131.110.4
Connecting to www.uca.edu.sv (www.uca.edu.sv)|201.131.110.4|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 274 [text/html]
Saving to: ‘/dev/null’

     0K                                                       100%  606M=0s

2020-02-25 22:13:22 (606 Mb/s) - ‘/dev/null’ saved [274/274]

--2020-02-25 22:13:22--  http://www.uca.edu.sv/-1DUgTd%0D
Resolving www.uca.edu.sv (www.uca.edu.sv)... 201.131.110.4
Connecting to www.uca.edu.sv (www.uca.edu.sv)|201.131.110.4|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 274 [text/html]
Saving to: ‘/dev/null’

     0K                                                       100%  718M=0s

2020-02-25 22:13:22 (718 Mb/s) - ‘/dev/null’ saved [274/274]

