--2020-03-02 03:27:29--  http://www.uma.edu.sv/image/pdf/diplomado.pdf
Resolving www.uma.edu.sv (www.uma.edu.sv)... 200.30.138.51
Connecting to www.uma.edu.sv (www.uma.edu.sv)|200.30.138.51|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 524227 (512K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  9% 1.55M 2s
    50K .......... .......... .......... .......... .......... 19% 1.74M 2s
   100K .......... .......... .......... .......... .......... 29% 3.17M 2s
   150K .......... .......... .......... .......... .......... 39% 11.5M 1s
   200K .......... .......... .......... .......... .......... 48% 4.08M 1s
   250K .......... .......... .......... .......... .......... 58% 12.6M 1s
   300K .......... .......... .......... .......... .......... 68% 4.08M 0s
   350K .......... .......... .......... .......... .......... 78% 14.9M 0s
   400K .......... .......... .......... .......... .......... 87% 94.5M 0s
   450K .......... .......... .......... .......... .......... 97% 4.03M 0s
   500K .......... .                                          100%  122M=1.0s

2020-03-02 03:27:31 (4.06 Mb/s) - ‘/dev/null’ saved [524227/524227]

