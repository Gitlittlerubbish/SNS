--2020-03-02 03:27:07--  http://www.insaforp.org.sv/siab/publicaciones/insaper36.pdf
Resolving www.insaforp.org.sv (www.insaforp.org.sv)... 66.198.240.17
Connecting to www.insaforp.org.sv (www.insaforp.org.sv)|66.198.240.17|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 81226 (79K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 63% 2.07M 0s
    50K .......... .......... .........                       100% 2.42M=0.3s

2020-03-02 03:27:07 (2.19 Mb/s) - ‘/dev/null’ saved [81226/81226]

