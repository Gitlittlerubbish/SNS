--2020-03-02 03:27:07--  http://libroslibres.uls.edu.sv/politica/militares_junto_al_pueblo.pdf
Resolving libroslibres.uls.edu.sv (libroslibres.uls.edu.sv)... 72.249.68.209
Connecting to libroslibres.uls.edu.sv (libroslibres.uls.edu.sv)|72.249.68.209|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 871306 (851K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  5% 1.87M 4s
    50K .......... .......... .......... .......... .......... 11% 3.69M 2s
   100K .......... .......... .......... .......... .......... 17% 30.9M 2s
   150K .......... .......... .......... .......... .......... 23% 4.45M 1s
   200K .......... .......... .......... .......... .......... 29% 51.5M 1s
   250K .......... .......... .......... .......... .......... 35% 26.7M 1s
   300K .......... .......... .......... .......... .......... 41% 4.48M 1s
   350K .......... .......... .......... .......... .......... 47% 67.5M 1s
   400K .......... .......... .......... .......... .......... 52%  113M 0s
   450K .......... .......... .......... .......... .......... 58% 32.8M 0s
   500K .......... .......... .......... .......... .......... 64% 4.33M 0s
   550K .......... .......... .......... .......... .......... 70%  140M 0s
   600K .......... .......... .......... .......... .......... 76% 85.2M 0s
   650K .......... .......... .......... .......... .......... 82% 81.5M 0s
   700K .......... .......... .......... .......... .......... 88% 55.2M 0s
   750K .......... .......... .......... .......... .......... 94% 4.26M 0s
   800K .......... .......... .......... .......... .......... 99%  339M 0s
   850K                                                       100%  145K=0.8s

2020-03-02 03:27:09 (8.89 Mb/s) - ‘/dev/null’ saved [871306/871306]

