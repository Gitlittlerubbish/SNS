--2020-02-25 22:13:40--  https://www.mh.gob.sv/downloads/pdf/PMHDC8306.pdf%0D
Resolving www.mh.gob.sv (www.mh.gob.sv)... 190.5.131.13, 190.57.24.24
Connecting to www.mh.gob.sv (www.mh.gob.sv)|190.5.131.13|:443... connected.
HTTP request sent, awaiting response... 302 Found
Location: https://www.mh.gob.sv/pmh/es/ [following]
--2020-02-25 22:13:41--  https://www.mh.gob.sv/pmh/es/
Reusing existing connection to www.mh.gob.sv:443.
HTTP request sent, awaiting response... 200 OK
Length: 57085 (56K) [text/html]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 89% 3.04M 0s
    50K .....                                                 100%  450M=0.1s

2020-02-25 22:13:41 (3.39 Mb/s) - ‘/dev/null’ saved [57085/57085]

--2020-02-25 22:13:41--  https://www.mh.gob.sv/downloads/pdf/PMHDC8306.pdf%0D
Resolving www.mh.gob.sv (www.mh.gob.sv)... 190.5.131.13, 190.57.24.24
Connecting to www.mh.gob.sv (www.mh.gob.sv)|190.5.131.13|:443... connected.
HTTP request sent, awaiting response... 302 Found
Location: https://www.mh.gob.sv/pmh/es/ [following]
--2020-02-25 22:13:41--  https://www.mh.gob.sv/pmh/es/
Reusing existing connection to www.mh.gob.sv:443.
HTTP request sent, awaiting response... 200 OK
Length: 57085 (56K) [text/html]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 89% 1.54M 0s
    50K .....                                                 100% 72.0M=0.3s

2020-02-25 22:13:42 (1.72 Mb/s) - ‘/dev/null’ saved [57085/57085]

--2020-02-25 22:14:10--  https://www.mh.gob.sv/downloads/pdf/PMHDC8306.pdf%0D
Resolving www.mh.gob.sv (www.mh.gob.sv)... 190.57.24.24, 190.5.131.13
Connecting to www.mh.gob.sv (www.mh.gob.sv)|190.57.24.24|:443... connected.
HTTP request sent, awaiting response... 302 Found
Location: https://www.mh.gob.sv/pmh/es/ [following]
--2020-02-25 22:14:10--  https://www.mh.gob.sv/pmh/es/
Reusing existing connection to www.mh.gob.sv:443.
HTTP request sent, awaiting response... 200 OK
Length: 57085 (56K) [text/html]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 89% 2.97M 0s
    50K .....                                                 100% 1.52G=0.1s

2020-02-25 22:14:10 (3.31 Mb/s) - ‘/dev/null’ saved [57085/57085]

--2020-02-25 22:14:10--  https://www.mh.gob.sv/downloads/pdf/PMHDC8306.pdf%0D
Resolving www.mh.gob.sv (www.mh.gob.sv)... 190.5.131.13, 190.57.24.24
Connecting to www.mh.gob.sv (www.mh.gob.sv)|190.5.131.13|:443... connected.
HTTP request sent, awaiting response... 302 Found
Location: https://www.mh.gob.sv/pmh/es/ [following]
--2020-02-25 22:14:11--  https://www.mh.gob.sv/pmh/es/
Reusing existing connection to www.mh.gob.sv:443.
HTTP request sent, awaiting response... 200 OK
Length: 57085 (56K) [text/html]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 89% 3.13M 0s
    50K .....                                                 100%  322M=0.1s

2020-02-25 22:14:11 (3.48 Mb/s) - ‘/dev/null’ saved [57085/57085]

