--2020-02-25 22:13:56--  http://www.insaforp.org.sv/siab/publicaciones/insaper36.pdf%0D
Resolving www.insaforp.org.sv (www.insaforp.org.sv)... 66.198.240.17
Connecting to www.insaforp.org.sv (www.insaforp.org.sv)|66.198.240.17|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:57 ERROR 404: Not Found.

--2020-02-25 22:14:23--  http://www.insaforp.org.sv/siab/publicaciones/insaper36.pdf%0D
Resolving www.insaforp.org.sv (www.insaforp.org.sv)... 66.198.240.17
Connecting to www.insaforp.org.sv (www.insaforp.org.sv)|66.198.240.17|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:23 ERROR 404: Not Found.

