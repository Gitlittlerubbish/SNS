--2020-02-25 22:12:55--  http://www.snet.gob.sv/Geologia/DeslavePicacho.pdf%0D
Resolving www.snet.gob.sv (www.snet.gob.sv)... 190.5.148.229, 170.0.177.4
Connecting to www.snet.gob.sv (www.snet.gob.sv)|190.5.148.229|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:12:55 ERROR 404: Not Found.

--2020-02-25 22:13:30--  http://www.snet.gob.sv/Geologia/DeslavePicacho.pdf%0D
Resolving www.snet.gob.sv (www.snet.gob.sv)... 170.0.177.4, 190.5.148.229
Connecting to www.snet.gob.sv (www.snet.gob.sv)|170.0.177.4|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:31 ERROR 404: Not Found.

