--2020-03-02 03:27:18--  http://tecnobodega.com.sv/images/Productos/20170620311528_V7S36LA.pdf
Resolving tecnobodega.com.sv (tecnobodega.com.sv)... 168.243.50.98
Connecting to tecnobodega.com.sv (tecnobodega.com.sv)|168.243.50.98|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 525409 (513K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  9%  968K 4s
    50K .......... .......... .......... .......... .......... 19% 2.97M 2s
   100K .......... .......... .......... .......... .......... 29% 71.5M 1s
   150K .......... .......... .......... .......... .......... 38% 1.47M 1s
   200K .......... .......... .......... .......... .......... 48%  419M 1s
   250K .......... .......... .......... .......... .......... 58% 2.91M 1s
   300K .......... .......... .......... .......... .......... 68% 1.46M 1s
   350K .......... .......... .......... .......... .......... 77% 3.20M 0s
   400K .......... .......... .......... .......... .......... 87% 2.72M 0s
   450K .......... .......... .......... .......... .......... 97% 2.91M 0s
   500K .......... ...                                        100%  797K=1.8s

2020-03-02 03:27:20 (2.31 Mb/s) - ‘/dev/null’ saved [525409/525409]

