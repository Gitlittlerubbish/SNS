--2020-03-02 03:24:32--  http://www.ute.gob.sv/publicaciones/0002.pdf
Resolving www.ute.gob.sv (www.ute.gob.sv)... 190.86.186.18
Connecting to www.ute.gob.sv (www.ute.gob.sv)|190.86.186.18|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 7951372 (7.6M) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  0% 1.33M 48s
    50K .......... .......... .......... .......... ..........  1% 2.38M 37s
   100K .......... .......... .......... .......... ..........  1% 2.47M 33s
   150K .......... .......... .......... .......... ..........  2% 2.47M 31s
   200K .......... .......... .......... .......... ..........  3% 2.46M 29s
   250K .......... .......... .......... .......... ..........  3% 2.47M 28s
   300K .......... .......... .......... .......... ..........  4% 2.45M 28s
   350K .......... .......... .......... .......... ..........  5% 2.48M 27s
   400K .......... .......... .......... .......... ..........  5% 2.39M 27s
   450K .......... .......... .......... .......... ..........  6% 2.48M 26s
   500K .......... .......... .......... .......... ..........  7% 2.45M 26s
   550K .......... .......... .......... .......... ..........  7% 2.46M 26s
   600K .......... .......... .......... .......... ..........  8% 2.44M 25s
   650K .......... .......... .......... .......... ..........  9% 2.46M 25s
   700K .......... .......... .......... .......... ..........  9% 2.40M 25s
   750K .......... .......... .......... .......... .......... 10% 2.45M 25s
   800K .......... .......... .......... .......... .......... 10% 2.46M 24s
   850K .......... .......... .......... .......... .......... 11% 2.46M 24s
   900K .......... .......... .......... .......... .......... 12% 2.47M 24s
   950K .......... .......... .......... .......... .......... 12% 2.40M 24s
  1000K .......... .......... .......... .......... .......... 13% 2.44M 23s
  1050K .......... .......... .......... .......... .......... 14% 2.47M 23s
  1100K .......... .......... .......... .......... .......... 14% 2.48M 23s
  1150K .......... .......... .......... .......... .......... 15% 2.43M 23s
  1200K .......... .......... .......... .......... .......... 16% 2.47M 23s
  1250K .......... .......... .......... .......... .......... 16% 2.43M 22s
  1300K .......... .......... .......... .......... .......... 17% 2.39M 22s
  1350K .......... .......... .......... .......... .......... 18% 2.48M 22s
  1400K .......... .......... .......... .......... .......... 18% 2.44M 22s
  1450K .......... .......... .......... .......... .......... 19% 2.46M 22s
  1500K .......... .......... .......... .......... .......... 19% 2.45M 21s
  1550K .......... .......... .......... .......... .......... 20% 2.46M 21s
  1600K .......... .......... .......... .......... .......... 21% 2.40M 21s
  1650K .......... .......... .......... .......... .......... 21% 2.44M 21s
  1700K .......... .......... .......... .......... .......... 22% 2.47M 21s
  1750K .......... .......... .......... .......... .......... 23% 2.44M 20s
  1800K .......... .......... .......... .......... .......... 23% 2.47M 20s
  1850K .......... .......... .......... .......... .......... 24% 2.46M 20s
  1900K .......... .......... .......... .......... .......... 25% 2.42M 20s
  1950K .......... .......... .......... .......... .......... 25% 2.41M 20s
  2000K .......... .......... .......... .......... .......... 26% 2.46M 20s
  2050K .......... .......... .......... .......... .......... 27% 2.46M 19s
  2100K .......... .......... .......... .......... .......... 27% 2.46M 19s
  2150K .......... .......... .......... .......... .......... 28% 2.45M 19s
  2200K .......... .......... .......... .......... .......... 28% 2.39M 19s
  2250K .......... .......... .......... .......... .......... 29% 2.49M 19s
  2300K .......... .......... .......... .......... .......... 30% 2.44M 18s
  2350K .......... .......... .......... .......... .......... 30% 2.44M 18s
  2400K .......... .......... .......... .......... .......... 31% 2.45M 18s
  2450K .......... .......... .......... .......... .......... 32% 2.45M 18s
  2500K .......... .......... .......... .......... .......... 32% 2.48M 18s
  2550K .......... .......... .......... .......... .......... 33% 2.45M 18s
  2600K .......... .......... .......... .......... .......... 34% 2.38M 17s
  2650K .......... .......... .......... .......... .......... 34% 2.43M 17s
  2700K .......... .......... .......... .......... .......... 35% 2.49M 17s
  2750K .......... .......... .......... .......... .......... 36% 2.45M 17s
  2800K .......... .......... .......... .......... .......... 36% 2.42M 17s
  2850K .......... .......... .......... .......... .......... 37% 2.41M 17s
  2900K .......... .......... .......... .......... .......... 37% 2.44M 16s
  2950K .......... .......... .......... .......... .......... 38% 2.48M 16s
  3000K .......... .......... .......... .......... .......... 39% 2.44M 16s
  3050K .......... .......... .......... .......... .......... 39% 2.45M 16s
  3100K .......... .......... .......... .......... .......... 40% 2.46M 16s
  3150K .......... .......... .......... .......... .......... 41% 2.46M 15s
  3200K .......... .......... .......... .......... .......... 41% 2.45M 15s
  3250K .......... .......... .......... .......... .......... 42% 2.39M 15s
  3300K .......... .......... .......... .......... .......... 43% 2.45M 15s
  3350K .......... .......... .......... .......... .......... 43% 2.46M 15s
  3400K .......... .......... .......... .......... .......... 44% 2.48M 15s
  3450K .......... .......... .......... .......... .......... 45% 2.43M 14s
  3500K .......... .......... .......... .......... .......... 45% 2.42M 14s
  3550K .......... .......... .......... .......... .......... 46% 2.44M 14s
  3600K .......... .......... .......... .......... .......... 47% 2.47M 14s
  3650K .......... .......... .......... .......... .......... 47% 2.47M 14s
  3700K .......... .......... .......... .......... .......... 48% 2.44M 14s
  3750K .......... .......... .......... .......... .......... 48% 2.47M 13s
  3800K .......... .......... .......... .......... .......... 49% 2.41M 13s
  3850K .......... .......... .......... .......... .......... 50% 2.46M 13s
  3900K .......... .......... .......... .......... .......... 50% 2.46M 13s
  3950K .......... .......... .......... .......... .......... 51% 2.44M 13s
  4000K .......... .......... .......... .......... .......... 52% 2.47M 13s
  4050K .......... .......... .......... .......... .......... 52% 2.46M 12s
  4100K .......... .......... .......... .......... .......... 53% 2.47M 12s
  4150K .......... .......... .......... .......... .......... 54% 2.46M 12s
  4200K .......... .......... .......... .......... .......... 54% 2.38M 12s
  4250K .......... .......... .......... .......... .......... 55% 2.46M 12s
  4300K .......... .......... .......... .......... .......... 56% 2.47M 12s
  4350K .......... .......... .......... .......... .......... 56% 2.47M 11s
  4400K .......... .......... .......... .......... .......... 57% 2.45M 11s
  4450K .......... .......... .......... .......... .......... 57% 2.39M 11s
  4500K .......... .......... .......... .......... .......... 58% 2.47M 11s
  4550K .......... .......... .......... .......... .......... 59% 2.46M 11s
  4600K .......... .......... .......... .......... .......... 59% 2.46M 11s
  4650K .......... .......... .......... .......... .......... 60% 2.47M 10s
  4700K .......... .......... .......... .......... .......... 61% 2.46M 10s
  4750K .......... .......... .......... .......... .......... 61% 2.45M 10s
  4800K .......... .......... .......... .......... .......... 62% 2.47M 10s
  4850K .......... .......... .......... .......... .......... 63% 2.37M 10s
  4900K .......... .......... .......... .......... .......... 63% 2.49M 10s
  4950K .......... .......... .......... .......... .......... 64% 2.47M 9s
  5000K .......... .......... .......... .......... .......... 65% 2.46M 9s
  5050K .......... .......... .......... .......... .......... 65% 2.45M 9s
  5100K .......... .......... .......... .......... .......... 66% 2.40M 9s
  5150K .......... .......... .......... .......... .......... 66% 2.46M 9s
  5200K .......... .......... .......... .......... .......... 67% 2.45M 8s
  5250K .......... .......... .......... .......... .......... 68% 2.46M 8s
  5300K .......... .......... .......... .......... .......... 68% 2.47M 8s
  5350K .......... .......... .......... .......... .......... 69% 2.45M 8s
  5400K .......... .......... .......... .......... .......... 70% 2.45M 8s
  5450K .......... .......... .......... .......... .......... 70% 2.49M 8s
  5500K .......... .......... .......... .......... .......... 71% 2.38M 7s
  5550K .......... .......... .......... .......... .......... 72% 2.46M 7s
  5600K .......... .......... .......... .......... .......... 72% 2.46M 7s
  5650K .......... .......... .......... .......... .......... 73% 2.46M 7s
  5700K .......... .......... .......... .......... .......... 74% 2.47M 7s
  5750K .......... .......... .......... .......... .......... 74% 2.39M 7s
  5800K .......... .......... .......... .......... .......... 75% 2.46M 6s
  5850K .......... .......... .......... .......... .......... 75% 2.45M 6s
  5900K .......... .......... .......... .......... .......... 76% 2.48M 6s
  5950K .......... .......... .......... .......... .......... 77% 2.46M 6s
  6000K .......... .......... .......... .......... .......... 77% 2.46M 6s
  6050K .......... .......... .......... .......... .......... 78% 2.46M 6s
  6100K .......... .......... .......... .......... .......... 79% 2.38M 5s
  6150K .......... .......... .......... .......... .......... 79% 2.47M 5s
  6200K .......... .......... .......... .......... .......... 80% 2.47M 5s
  6250K .......... .......... .......... .......... .......... 81% 2.46M 5s
  6300K .......... .......... .......... .......... .......... 81% 2.47M 5s
  6350K .......... .......... .......... .......... .......... 82% 2.47M 5s
  6400K .......... .......... .......... .......... .......... 83% 2.39M 4s
  6450K .......... .......... .......... .......... .......... 83% 2.44M 4s
  6500K .......... .......... .......... .......... .......... 84% 2.47M 4s
  6550K .......... .......... .......... .......... .......... 84% 2.45M 4s
  6600K .......... .......... .......... .......... .......... 85% 2.46M 4s
  6650K .......... .......... .......... .......... .......... 86% 2.48M 4s
  6700K .......... .......... .......... .......... .......... 86% 2.46M 3s
  6750K .......... .......... .......... .......... .......... 87% 2.40M 3s
  6800K .......... .......... .......... .......... .......... 88% 2.46M 3s
  6850K .......... .......... .......... .......... .......... 88% 2.46M 3s
  6900K .......... .......... .......... .......... .......... 89% 2.48M 3s
  6950K .......... .......... .......... .......... .......... 90% 2.44M 3s
  7000K .......... .......... .......... .......... .......... 90% 2.41M 2s
  7050K .......... .......... .......... .......... .......... 91% 2.46M 2s
  7100K .......... .......... .......... .......... .......... 92% 2.45M 2s
  7150K .......... .......... .......... .......... .......... 92% 2.48M 2s
  7200K .......... .......... .......... .......... .......... 93% 2.43M 2s
  7250K .......... .......... .......... .......... .......... 94% 2.48M 2s
  7300K .......... .......... .......... .......... .......... 94% 2.48M 1s
  7350K .......... .......... .......... .......... .......... 95% 2.35M 1s
  7400K .......... .......... .......... .......... .......... 95% 2.49M 1s
  7450K .......... .......... .......... .......... .......... 96% 2.47M 1s
  7500K .......... .......... .......... .......... .......... 97% 2.47M 1s
  7550K .......... .......... .......... .......... .......... 97% 2.46M 1s
  7600K .......... .......... .......... .......... .......... 98% 2.45M 0s
  7650K .......... .......... .......... .......... .......... 99% 2.46M 0s
  7700K .......... .......... .......... .......... .......... 99% 2.41M 0s
  7750K .......... .....                                      100% 1.11M=26s

2020-03-02 03:24:59 (2.43 Mb/s) - ‘/dev/null’ saved [7951372/7951372]

