--2020-03-02 03:26:23--  http://www.ugb.edu.sv/images/pdf/modeloeducativougb.pdf
Resolving www.ugb.edu.sv (www.ugb.edu.sv)... 190.86.248.10
Connecting to www.ugb.edu.sv (www.ugb.edu.sv)|190.86.248.10|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 1154724 (1.1M) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  4%  233K 38s
    50K .......... .......... .......... .......... ..........  8%  182K 41s
   100K .......... .......... .......... .......... .......... 13%  171K 42s
   150K .......... .......... .......... .......... .......... 17%  181K 40s
   200K .......... .......... .......... .......... .......... 22%  165K 39s
   250K .......... .......... .......... .......... .......... 26%  234K 36s
   300K .......... .......... .......... .......... .......... 31%  194K 33s
   350K .......... .......... .......... .......... .......... 35%  196K 31s
   400K .......... .......... .......... .......... .......... 39%  169K 29s
   450K .......... .......... .......... .......... .......... 44%  207K 27s
   500K .......... .......... .......... .......... .......... 48%  217K 25s
   550K .......... .......... .......... .......... .......... 53%  285K 22s
   600K .......... .......... .......... .......... .......... 57%  202K 20s
   650K .......... .......... .......... .......... .......... 62%  193K 18s
   700K .......... .......... .......... .......... .......... 66%  232K 15s
   750K .......... .......... .......... .......... .......... 70%  226K 13s
   800K .......... .......... .......... .......... .......... 75%  327K 11s
   850K .......... .......... .......... .......... .......... 79%  288K 9s
   900K .......... .......... .......... .......... .......... 84%  251K 7s
   950K .......... .......... .......... .......... .......... 88%  238K 5s
  1000K .......... .......... .......... .......... .......... 93%  221K 3s
  1050K .......... .......... .......... .......... .......... 97%  233K 1s
  1100K .......... .......... .......                         100%  290K=43s

2020-03-02 03:27:07 (215 Kb/s) - ‘/dev/null’ saved [1154724/1154724]

