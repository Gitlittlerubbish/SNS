--2020-03-02 03:25:39--  http://www.evivienda.gob.sv/Lotificaciones/Documentos/INSTRUCTIVO_SIL.pdf
Resolving www.evivienda.gob.sv (www.evivienda.gob.sv)... 200.31.181.149
Connecting to www.evivienda.gob.sv (www.evivienda.gob.sv)|200.31.181.149|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 1488648 (1.4M) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  3% 1.02M 11s
    50K .......... .......... .......... .......... ..........  6% 1.08M 11s
   100K .......... .......... .......... .......... .......... 10%  912K 11s
   150K .......... .......... .......... .......... .......... 13% 1.23M 10s
   200K .......... .......... .......... .......... .......... 17%  849K 10s
   250K .......... .......... .......... .......... .......... 20% 1.02M 9s
   300K .......... .......... .......... .......... .......... 24%  912K 9s
   350K .......... .......... .......... .......... .......... 27% 1.02M 9s
   400K .......... .......... .......... .......... .......... 30% 1.08M 8s
   450K .......... .......... .......... .......... .......... 34%  962K 8s
   500K .......... .......... .......... .......... .......... 37% 1.11M 7s
   550K .......... .......... .......... .......... .......... 41% 1.05M 7s
   600K .......... .......... .......... .......... .......... 44%  790K 7s
   650K .......... .......... .......... .......... .......... 48% 1.19M 6s
   700K .......... .......... .......... .......... .......... 51%  826K 6s
   750K .......... .......... .......... .......... .......... 55% 1.56M 5s
   800K .......... .......... .......... .......... .......... 58%  806K 5s
   850K .......... .......... .......... .......... .......... 61%  939K 5s
   900K .......... .......... .......... .......... .......... 65%  895K 4s
   950K .......... .......... .......... .......... .......... 68% 1.18M 4s
  1000K .......... .......... .......... .......... .......... 72% 1.08M 3s
  1050K .......... .......... .......... .......... .......... 75% 1.08M 3s
  1100K .......... .......... .......... .......... .......... 79%  890K 2s
  1150K .......... .......... .......... .......... .......... 82%  867K 2s
  1200K .......... .......... .......... .......... .......... 85% 1.12M 2s
  1250K .......... .......... .......... .......... .......... 89%  890K 1s
  1300K .......... .......... .......... .......... .......... 92% 1.23M 1s
  1350K .......... .......... .......... .......... .......... 96% 1.12M 0s
  1400K .......... .......... .......... .......... .......... 99%  790K 0s
  1450K ...                                                   100%  327K=12s

2020-03-02 03:25:52 (987 Kb/s) - ‘/dev/null’ saved [1488648/1488648]

