--2020-03-02 03:25:38--  http://puntosdeventa.com.sv/manuales/47/DS000003_1515L.pdf
Resolving puntosdeventa.com.sv (puntosdeventa.com.sv)... 67.227.226.242
Connecting to puntosdeventa.com.sv (puntosdeventa.com.sv)|67.227.226.242|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 320849 (313K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 15% 2.02M 1s
    50K .......... .......... .......... .......... .......... 31% 4.01M 1s
   100K .......... .......... .......... .......... .......... 47% 4.03M 0s
   150K .......... .......... .......... .......... .......... 63% 4.10M 0s
   200K .......... .......... .......... .......... .......... 79%  198M 0s
   250K .......... .......... .......... .......... .......... 95% 4.18M 0s
   300K .......... ...                                        100%  691M=0.6s

2020-03-02 03:25:39 (4.23 Mb/s) - ‘/dev/null’ saved [320849/320849]

