--2020-02-25 22:12:46--  http://appm.aduana.gob.sv/sacelectronico/NOTAS%2520EXPLICATIVAS.pdf%0D
Resolving appm.aduana.gob.sv (appm.aduana.gob.sv)... 190.5.131.16, 190.57.24.28
Connecting to appm.aduana.gob.sv (appm.aduana.gob.sv)|190.5.131.16|:80... connected.
HTTP request sent, awaiting response... 400 Bad Request
2020-02-25 22:12:47 ERROR 400: Bad Request.

--2020-02-25 22:13:24--  http://appm.aduana.gob.sv/sacelectronico/NOTAS%2520EXPLICATIVAS.pdf%0D
Resolving appm.aduana.gob.sv (appm.aduana.gob.sv)... 190.5.131.16, 190.57.24.28
Connecting to appm.aduana.gob.sv (appm.aduana.gob.sv)|190.5.131.16|:80... connected.
HTTP request sent, awaiting response... 400 Bad Request
2020-02-25 22:13:25 ERROR 400: Bad Request.

