--2020-02-25 22:12:27--  http://biblioteca.ues.edu.sv/revistas/10800099.pdf%0D
Resolving biblioteca.ues.edu.sv (biblioteca.ues.edu.sv)... 168.232.48.132
Connecting to biblioteca.ues.edu.sv (biblioteca.ues.edu.sv)|168.232.48.132|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:12:31 ERROR 404: Not Found.

--2020-02-25 22:12:31--  http://biblioteca.ues.edu.sv/revistas/10800057E1.pdf%0D
Resolving biblioteca.ues.edu.sv (biblioteca.ues.edu.sv)... 168.232.48.132
Connecting to biblioteca.ues.edu.sv (biblioteca.ues.edu.sv)|168.232.48.132|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:12:31 ERROR 404: Not Found.

--2020-02-25 22:13:15--  http://biblioteca.ues.edu.sv/revistas/10800099.pdf%0D
Resolving biblioteca.ues.edu.sv (biblioteca.ues.edu.sv)... 168.232.48.132
Connecting to biblioteca.ues.edu.sv (biblioteca.ues.edu.sv)|168.232.48.132|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:15 ERROR 404: Not Found.

--2020-02-25 22:13:15--  http://biblioteca.ues.edu.sv/revistas/10800057E1.pdf%0D
Resolving biblioteca.ues.edu.sv (biblioteca.ues.edu.sv)... 168.232.48.132
Connecting to biblioteca.ues.edu.sv (biblioteca.ues.edu.sv)|168.232.48.132|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:15 ERROR 404: Not Found.

