--2020-02-25 22:12:49--  http://www.brasil.org.sv/Paginas/Orientacao.pdf%0D
Resolving www.brasil.org.sv (www.brasil.org.sv)... failed: Name or service not known.
wget: unable to resolve host address ‘www.brasil.org.sv’
--2020-02-25 22:13:26--  http://www.brasil.org.sv/Paginas/Orientacao.pdf%0D
Resolving www.brasil.org.sv (www.brasil.org.sv)... failed: Name or service not known.
wget: unable to resolve host address ‘www.brasil.org.sv’
