--2020-02-25 22:13:54--  https://ui.usonsonate.edu.sv/papers/DIRECTORES_EXITOSOS.pdf%0D
Resolving ui.usonsonate.edu.sv (ui.usonsonate.edu.sv)... 66.113.161.172
Connecting to ui.usonsonate.edu.sv (ui.usonsonate.edu.sv)|66.113.161.172|:443... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:54 ERROR 404: Not Found.

--2020-02-25 22:14:20--  https://ui.usonsonate.edu.sv/papers/DIRECTORES_EXITOSOS.pdf%0D
Resolving ui.usonsonate.edu.sv (ui.usonsonate.edu.sv)... 66.113.161.172
Connecting to ui.usonsonate.edu.sv (ui.usonsonate.edu.sv)|66.113.161.172|:443... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:21 ERROR 404: Not Found.

