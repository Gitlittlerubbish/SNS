--2020-03-02 03:24:13--  http://www.amway.com.sv/downloads/Catalogo_Nutrilite_2015.pdf
Resolving www.amway.com.sv (www.amway.com.sv)... 92.123.196.133
Connecting to www.amway.com.sv (www.amway.com.sv)|92.123.196.133|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 23622382 (23M) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  0% 60.4M 3s
    50K .......... .......... .......... .......... ..........  0% 71.7M 3s
   100K .......... .......... .......... .......... ..........  0%  128M 2s
   150K .......... .......... .......... .......... ..........  0%  109M 2s
   200K .......... .......... .......... .......... ..........  1%  505M 2s
   250K .......... .......... .......... .......... ..........  1% 69.0M 2s
   300K .......... .......... .......... .......... ..........  1%  134M 2s
   350K .......... .......... .......... .......... ..........  1%  406M 2s
   400K .......... .......... .......... .......... ..........  1%  193M 2s
   450K .......... .......... .......... .......... ..........  2%  235M 2s
   500K .......... .......... .......... .......... ..........  2% 98.9M 2s
   550K .......... .......... .......... .......... ..........  2%  143M 2s
   600K .......... .......... .......... .......... ..........  2% 1.70G 1s
   650K .......... .......... .......... .......... ..........  3%  217M 1s
   700K .......... .......... .......... .......... ..........  3%  474M 1s
   750K .......... .......... .......... .......... ..........  3%  415M 1s
   800K .......... .......... .......... .......... ..........  3%  208M 1s
   850K .......... .......... .......... .......... ..........  3%  443M 1s
   900K .......... .......... .......... .......... ..........  4% 89.4M 1s
   950K .......... .......... .......... .......... ..........  4%  206M 1s
  1000K .......... .......... .......... .......... ..........  4%  388M 1s
  1050K .......... .......... .......... .......... ..........  4%  355M 1s
  1100K .......... .......... .......... .......... ..........  4%  326M 1s
  1150K .......... .......... .......... .......... ..........  5%  239M 1s
  1200K .......... .......... .......... .......... ..........  5% 63.1M 1s
  1250K .......... .......... .......... .......... ..........  5%  306M 1s
  1300K .......... .......... .......... .......... ..........  5%  331M 1s
  1350K .......... .......... .......... .......... ..........  6%  275M 1s
  1400K .......... .......... .......... .......... ..........  6%  187M 1s
  1450K .......... .......... .......... .......... ..........  6%  237M 1s
  1500K .......... .......... .......... .......... ..........  6% 24.3M 1s
  1550K .......... .......... .......... .......... ..........  6%  423M 1s
  1600K .......... .......... .......... .......... ..........  7%  502M 1s
  1650K .......... .......... .......... .......... ..........  7%  256M 1s
  1700K .......... .......... .......... .......... ..........  7%  363M 1s
  1750K .......... .......... .......... .......... ..........  7% 99.5M 1s
  1800K .......... .......... .......... .......... ..........  8%  746M 1s
  1850K .......... .......... .......... .......... ..........  8%  230M 1s
  1900K .......... .......... .......... .......... ..........  8% 89.4M 1s
  1950K .......... .......... .......... .......... ..........  8% 9.18M 2s
  2000K .......... .......... .......... .......... ..........  8% 1.97G 2s
  2050K .......... .......... .......... .......... ..........  9% 1.90G 2s
  2100K .......... .......... .......... .......... ..........  9% 2.11G 1s
  2150K .......... .......... .......... .......... ..........  9% 2.41G 1s
  2200K .......... .......... .......... .......... ..........  9% 2.38G 1s
  2250K .......... .......... .......... .......... ..........  9% 2.59G 1s
  2300K .......... .......... .......... .......... .......... 10%  160M 1s
  2350K .......... .......... .......... .......... .......... 10% 78.4M 1s
  2400K .......... .......... .......... .......... .......... 10% 12.1M 2s
  2450K .......... .......... .......... .......... .......... 10%  178M 2s
  2500K .......... .......... .......... .......... .......... 11%  506M 2s
  2550K .......... .......... .......... .......... .......... 11%  127M 2s
  2600K .......... .......... .......... .......... .......... 11% 19.7M 2s
  2650K .......... .......... .......... .......... .......... 11% 2.59G 2s
  2700K .......... .......... .......... .......... .......... 11% 2.95G 2s
  2750K .......... .......... .......... .......... .......... 12% 2.71G 2s
  2800K .......... .......... .......... .......... .......... 12% 3.15G 2s
  2850K .......... .......... .......... .......... .......... 12%  509M 2s
  2900K .......... .......... .......... .......... .......... 12%  130M 2s
  2950K .......... .......... .......... .......... .......... 13% 33.4M 2s
  3000K .......... .......... .......... .......... .......... 13% 65.6M 2s
  3050K .......... .......... .......... .......... .......... 13%  143M 2s
  3100K .......... .......... .......... .......... .......... 13%  283M 2s
  3150K .......... .......... .......... .......... .......... 13% 64.0M 2s
  3200K .......... .......... .......... .......... .......... 14% 67.3M 2s
  3250K .......... .......... .......... .......... .......... 14% 72.0M 2s
  3300K .......... .......... .......... .......... .......... 14% 65.0M 2s
  3350K .......... .......... .......... .......... .......... 14% 76.1M 2s
  3400K .......... .......... .......... .......... .......... 14% 51.2M 2s
  3450K .......... .......... .......... .......... .......... 15% 81.7M 2s
  3500K .......... .......... .......... .......... .......... 15% 80.1M 2s
  3550K .......... .......... .......... .......... .......... 15% 74.3M 2s
  3600K .......... .......... .......... .......... .......... 15% 63.2M 2s
  3650K .......... .......... .......... .......... .......... 16% 69.7M 2s
  3700K .......... .......... .......... .......... .......... 16% 65.3M 2s
  3750K .......... .......... .......... .......... .......... 16% 38.8M 2s
  3800K .......... .......... .......... .......... .......... 16%  181M 2s
  3850K .......... .......... .......... .......... .......... 16% 57.9M 2s
  3900K .......... .......... .......... .......... .......... 17% 60.0M 2s
  3950K .......... .......... .......... .......... .......... 17% 66.3M 2s
  4000K .......... .......... .......... .......... .......... 17% 82.6M 2s
  4050K .......... .......... .......... .......... .......... 17% 68.9M 2s
  4100K .......... .......... .......... .......... .......... 17%  103M 2s
  4150K .......... .......... .......... .......... .......... 18% 76.7M 2s
  4200K .......... .......... .......... .......... .......... 18% 79.5M 2s
  4250K .......... .......... .......... .......... .......... 18% 61.9M 2s
  4300K .......... .......... .......... .......... .......... 18% 61.4M 2s
  4350K .......... .......... .......... .......... .......... 19%  105M 2s
  4400K .......... .......... .......... .......... .......... 19% 55.1M 2s
  4450K .......... .......... .......... .......... .......... 19% 78.8M 2s
  4500K .......... .......... .......... .......... .......... 19% 66.2M 2s
  4550K .......... .......... .......... .......... .......... 19% 79.1M 2s
  4600K .......... .......... .......... .......... .......... 20% 74.1M 2s
  4650K .......... .......... .......... .......... .......... 20% 64.2M 2s
  4700K .......... .......... .......... .......... .......... 20% 55.2M 2s
  4750K .......... .......... .......... .......... .......... 20% 83.5M 2s
  4800K .......... .......... .......... .......... .......... 21% 70.4M 2s
  4850K .......... .......... .......... .......... .......... 21% 69.1M 2s
  4900K .......... .......... .......... .......... .......... 21% 75.7M 2s
  4950K .......... .......... .......... .......... .......... 21% 74.9M 2s
  5000K .......... .......... .......... .......... .......... 21% 63.2M 2s
  5050K .......... .......... .......... .......... .......... 22% 69.2M 2s
  5100K .......... .......... .......... .......... .......... 22% 72.5M 2s
  5150K .......... .......... .......... .......... .......... 22% 35.9M 2s
  5200K .......... .......... .......... .......... .......... 22% 83.1M 2s
  5250K .......... .......... .......... .......... .......... 22%  163M 2s
  5300K .......... .......... .......... .......... .......... 23% 62.3M 2s
  5350K .......... .......... .......... .......... .......... 23% 54.2M 2s
  5400K .......... .......... .......... .......... .......... 23%  100M 2s
  5450K .......... .......... .......... .......... .......... 23% 48.9M 2s
  5500K .......... .......... .......... .......... .......... 24%  104M 2s
  5550K .......... .......... .......... .......... .......... 24% 77.5M 2s
  5600K .......... .......... .......... .......... .......... 24% 87.3M 2s
  5650K .......... .......... .......... .......... .......... 24% 70.9M 2s
  5700K .......... .......... .......... .......... .......... 24% 60.1M 2s
  5750K .......... .......... .......... .......... .......... 25% 75.6M 2s
  5800K .......... .......... .......... .......... .......... 25% 67.7M 2s
  5850K .......... .......... .......... .......... .......... 25% 58.9M 2s
  5900K .......... .......... .......... .......... .......... 25% 79.1M 2s
  5950K .......... .......... .......... .......... .......... 26% 87.5M 2s
  6000K .......... .......... .......... .......... .......... 26% 76.9M 2s
  6050K .......... .......... .......... .......... .......... 26% 71.6M 2s
  6100K .......... .......... .......... .......... .......... 26% 60.6M 2s
  6150K .......... .......... .......... .......... .......... 26% 88.2M 2s
  6200K .......... .......... .......... .......... .......... 27% 72.4M 2s
  6250K .......... .......... .......... .......... .......... 27% 62.2M 2s
  6300K .......... .......... .......... .......... .......... 27% 93.4M 2s
  6350K .......... .......... .......... .......... .......... 27% 69.1M 2s
  6400K .......... .......... .......... .......... .......... 27% 79.0M 2s
  6450K .......... .......... .......... .......... .......... 28% 60.7M 2s
  6500K .......... .......... .......... .......... .......... 28% 84.9M 2s
  6550K .......... .......... .......... .......... .......... 28% 72.2M 2s
  6600K .......... .......... .......... .......... .......... 28% 72.2M 2s
  6650K .......... .......... .......... .......... .......... 29% 72.6M 2s
  6700K .......... .......... .......... .......... .......... 29% 74.4M 2s
  6750K .......... .......... .......... .......... .......... 29% 68.3M 2s
  6800K .......... .......... .......... .......... .......... 29% 29.0M 2s
  6850K .......... .......... .......... .......... .......... 29% 2.34G 2s
  6900K .......... .......... .......... .......... .......... 30%  160M 2s
  6950K .......... .......... .......... .......... .......... 30% 57.6M 2s
  7000K .......... .......... .......... .......... .......... 30% 66.7M 2s
  7050K .......... .......... .......... .......... .......... 30% 75.3M 2s
  7100K .......... .......... .......... .......... .......... 30% 77.4M 2s
  7150K .......... .......... .......... .......... .......... 31% 80.3M 2s
  7200K .......... .......... .......... .......... .......... 31% 81.3M 2s
  7250K .......... .......... .......... .......... .......... 31% 88.6M 2s
  7300K .......... .......... .......... .......... .......... 31% 69.3M 2s
  7350K .......... .......... .......... .......... .......... 32% 55.1M 2s
  7400K .......... .......... .......... .......... .......... 32%  109M 2s
  7450K .......... .......... .......... .......... .......... 32% 68.7M 2s
  7500K .......... .......... .......... .......... .......... 32% 83.2M 2s
  7550K .......... .......... .......... .......... .......... 32% 75.2M 2s
  7600K .......... .......... .......... .......... .......... 33% 74.3M 2s
  7650K .......... .......... .......... .......... .......... 33% 60.6M 2s
  7700K .......... .......... .......... .......... .......... 33% 77.7M 2s
  7750K .......... .......... .......... .......... .......... 33% 81.7M 2s
  7800K .......... .......... .......... .......... .......... 34% 75.5M 2s
  7850K .......... .......... .......... .......... .......... 34% 70.2M 2s
  7900K .......... .......... .......... .......... .......... 34% 74.1M 2s
  7950K .......... .......... .......... .......... .......... 34% 70.2M 2s
  8000K .......... .......... .......... .......... .......... 34% 73.7M 2s
  8050K .......... .......... .......... .......... .......... 35% 74.7M 2s
  8100K .......... .......... .......... .......... .......... 35% 42.4M 2s
  8150K .......... .......... .......... .......... .......... 35%  164M 2s
  8200K .......... .......... .......... .......... .......... 35% 62.5M 2s
  8250K .......... .......... .......... .......... .......... 35% 45.8M 2s
  8300K .......... .......... .......... .......... .......... 36% 58.4M 2s
  8350K .......... .......... .......... .......... .......... 36% 82.7M 2s
  8400K .......... .......... .......... .......... .......... 36% 67.5M 1s
  8450K .......... .......... .......... .......... .......... 36% 80.5M 1s
  8500K .......... .......... .......... .......... .......... 37% 80.6M 1s
  8550K .......... .......... .......... .......... .......... 37% 62.4M 1s
  8600K .......... .......... .......... .......... .......... 37% 11.1M 2s
  8650K .......... .......... .......... .......... .......... 37% 73.7M 2s
  8700K .......... .......... .......... .......... .......... 37% 90.1M 2s
  8750K .......... .......... .......... .......... .......... 38% 80.3M 2s
  8800K .......... .......... .......... .......... .......... 38% 94.0M 2s
  8850K .......... .......... .......... .......... .......... 38%  130M 2s
  8900K .......... .......... .......... .......... .......... 38% 84.6M 1s
  8950K .......... .......... .......... .......... .......... 39%  102M 1s
  9000K .......... .......... .......... .......... .......... 39%  103M 1s
  9050K .......... .......... .......... .......... .......... 39%  160M 1s
  9100K .......... .......... .......... .......... .......... 39% 93.7M 1s
  9150K .......... .......... .......... .......... .......... 39%  128M 1s
  9200K .......... .......... .......... .......... .......... 40%  108M 1s
  9250K .......... .......... .......... .......... .......... 40%  111M 1s
  9300K .......... .......... .......... .......... .......... 40%  115M 1s
  9350K .......... .......... .......... .......... .......... 40%  147M 1s
  9400K .......... .......... .......... .......... .......... 40% 98.9M 1s
  9450K .......... .......... .......... .......... .......... 41%  127M 1s
  9500K .......... .......... .......... .......... .......... 41% 5.02M 2s
  9550K .......... .......... .......... .......... .......... 41% 96.4M 2s
  9600K .......... .......... .......... .......... .......... 41%  121M 1s
  9650K .......... .......... .......... .......... .......... 42%  134M 1s
  9700K .......... .......... .......... .......... .......... 42%  137M 1s
  9750K .......... .......... .......... .......... .......... 42%  147M 1s
  9800K .......... .......... .......... .......... .......... 42% 94.4M 1s
  9850K .......... .......... .......... .......... .......... 42% 33.4M 1s
  9900K .......... .......... .......... .......... .......... 43%  109M 1s
  9950K .......... .......... .......... .......... .......... 43%  130M 1s
 10000K .......... .......... .......... .......... .......... 43%  102M 1s
 10050K .......... .......... .......... .......... .......... 43% 89.4M 1s
 10100K .......... .......... .......... .......... .......... 43% 77.8M 1s
 10150K .......... .......... .......... .......... .......... 44%  112M 1s
 10200K .......... .......... .......... .......... .......... 44% 74.9M 1s
 10250K .......... .......... .......... .......... .......... 44%  106M 1s
 10300K .......... .......... .......... .......... .......... 44%  127M 1s
 10350K .......... .......... .......... .......... .......... 45%  119M 1s
 10400K .......... .......... .......... .......... .......... 45% 91.0M 1s
 10450K .......... .......... .......... .......... .......... 45%  141M 1s
 10500K .......... .......... .......... .......... .......... 45% 79.8M 1s
 10550K .......... .......... .......... .......... .......... 45%  102M 1s
 10600K .......... .......... .......... .......... .......... 46%  146M 1s
 10650K .......... .......... .......... .......... .......... 46% 79.8M 1s
 10700K .......... .......... .......... .......... .......... 46%  137M 1s
 10750K .......... .......... .......... .......... .......... 46%  115M 1s
 10800K .......... .......... .......... .......... .......... 47%  181M 1s
 10850K .......... .......... .......... .......... .......... 47%  127M 1s
 10900K .......... .......... .......... .......... .......... 47%  128M 1s
 10950K .......... .......... .......... .......... .......... 47%  114M 1s
 11000K .......... .......... .......... .......... .......... 47%  183M 1s
 11050K .......... .......... .......... .......... .......... 48%  149M 1s
 11100K .......... .......... .......... .......... .......... 48%  128M 1s
 11150K .......... .......... .......... .......... .......... 48%  216M 1s
 11200K .......... .......... .......... .......... .......... 48%  127M 1s
 11250K .......... .......... .......... .......... .......... 48%  105M 1s
 11300K .......... .......... .......... .......... .......... 49%  145M 1s
 11350K .......... .......... .......... .......... .......... 49%  150M 1s
 11400K .......... .......... .......... .......... .......... 49%  117M 1s
 11450K .......... .......... .......... .......... .......... 49%  187M 1s
 11500K .......... .......... .......... .......... .......... 50%  155M 1s
 11550K .......... .......... .......... .......... .......... 50%  201M 1s
 11600K .......... .......... .......... .......... .......... 50%  159M 1s
 11650K .......... .......... .......... .......... .......... 50%  101M 1s
 11700K .......... .......... .......... .......... .......... 50% 77.4M 1s
 11750K .......... .......... .......... .......... .......... 51% 34.7M 1s
 11800K .......... .......... .......... .......... .......... 51%  525M 1s
 11850K .......... .......... .......... .......... .......... 51%  111M 1s
 11900K .......... .......... .......... .......... .......... 51% 70.7M 1s
 11950K .......... .......... .......... .......... .......... 52% 67.2M 1s
 12000K .......... .......... .......... .......... .......... 52% 77.4M 1s
 12050K .......... .......... .......... .......... .......... 52% 71.7M 1s
 12100K .......... .......... .......... .......... .......... 52% 75.6M 1s
 12150K .......... .......... .......... .......... .......... 52% 65.2M 1s
 12200K .......... .......... .......... .......... .......... 53% 88.0M 1s
 12250K .......... .......... .......... .......... .......... 53% 67.6M 1s
 12300K .......... .......... .......... .......... .......... 53% 83.5M 1s
 12350K .......... .......... .......... .......... .......... 53% 67.5M 1s
 12400K .......... .......... .......... .......... .......... 53% 74.0M 1s
 12450K .......... .......... .......... .......... .......... 54% 75.4M 1s
 12500K .......... .......... .......... .......... .......... 54% 54.7M 1s
 12550K .......... .......... .......... .......... .......... 54% 98.6M 1s
 12600K .......... .......... .......... .......... .......... 54% 76.4M 1s
 12650K .......... .......... .......... .......... .......... 55% 77.0M 1s
 12700K .......... .......... .......... .......... .......... 55% 68.7M 1s
 12750K .......... .......... .......... .......... .......... 55% 71.6M 1s
 12800K .......... .......... .......... .......... .......... 55% 82.3M 1s
 12850K .......... .......... .......... .......... .......... 55% 58.7M 1s
 12900K .......... .......... .......... .......... .......... 56% 92.6M 1s
 12950K .......... .......... .......... .......... .......... 56% 71.3M 1s
 13000K .......... .......... .......... .......... .......... 56% 76.8M 1s
 13050K .......... .......... .......... .......... .......... 56% 33.9M 1s
 13100K .......... .......... .......... .......... .......... 57% 3.20G 1s
 13150K .......... .......... .......... .......... .......... 57% 69.4M 1s
 13200K .......... .......... .......... .......... .......... 57% 95.3M 1s
 13250K .......... .......... .......... .......... .......... 57% 61.1M 1s
 13300K .......... .......... .......... .......... .......... 57% 77.3M 1s
 13350K .......... .......... .......... .......... .......... 58% 80.0M 1s
 13400K .......... .......... .......... .......... .......... 58% 62.4M 1s
 13450K .......... .......... .......... .......... .......... 58% 83.1M 1s
 13500K .......... .......... .......... .......... .......... 58% 73.6M 1s
 13550K .......... .......... .......... .......... .......... 58% 67.8M 1s
 13600K .......... .......... .......... .......... .......... 59% 85.5M 1s
 13650K .......... .......... .......... .......... .......... 59% 65.0M 1s
 13700K .......... .......... .......... .......... .......... 59% 69.6M 1s
 13750K .......... .......... .......... .......... .......... 59% 63.9M 1s
 13800K .......... .......... .......... .......... .......... 60% 82.5M 1s
 13850K .......... .......... .......... .......... .......... 60% 92.8M 1s
 13900K .......... .......... .......... .......... .......... 60% 68.3M 1s
 13950K .......... .......... .......... .......... .......... 60% 70.9M 1s
 14000K .......... .......... .......... .......... .......... 60% 77.4M 1s
 14050K .......... .......... .......... .......... .......... 61% 77.2M 1s
 14100K .......... .......... .......... .......... .......... 61% 74.4M 1s
 14150K .......... .......... .......... .......... .......... 61% 67.1M 1s
 14200K .......... .......... .......... .......... .......... 61% 66.6M 1s
 14250K .......... .......... .......... .......... .......... 61% 82.5M 1s
 14300K .......... .......... .......... .......... .......... 62% 77.1M 1s
 14350K .......... .......... .......... .......... .......... 62% 59.4M 1s
 14400K .......... .......... .......... .......... .......... 62% 77.6M 1s
 14450K .......... .......... .......... .......... .......... 62% 42.5M 1s
 14500K .......... .......... .......... .......... .......... 63%  433M 1s
 14550K .......... .......... .......... .......... .......... 63% 54.9M 1s
 14600K .......... .......... .......... .......... .......... 63% 88.9M 1s
 14650K .......... .......... .......... .......... .......... 63% 57.9M 1s
 14700K .......... .......... .......... .......... .......... 63% 68.7M 1s
 14750K .......... .......... .......... .......... .......... 64% 83.0M 1s
 14800K .......... .......... .......... .......... .......... 64% 77.6M 1s
 14850K .......... .......... .......... .......... .......... 64% 91.8M 1s
 14900K .......... .......... .......... .......... .......... 64% 75.7M 1s
 14950K .......... .......... .......... .......... .......... 65% 69.4M 1s
 15000K .......... .......... .......... .......... .......... 65% 76.7M 1s
 15050K .......... .......... .......... .......... .......... 65% 72.7M 1s
 15100K .......... .......... .......... .......... .......... 65% 75.7M 1s
 15150K .......... .......... .......... .......... .......... 65% 72.4M 1s
 15200K .......... .......... .......... .......... .......... 66% 68.2M 1s
 15250K .......... .......... .......... .......... .......... 66% 6.68M 1s
 15300K .......... .......... .......... .......... .......... 66% 83.5M 1s
 15350K .......... .......... .......... .......... .......... 66% 83.0M 1s
 15400K .......... .......... .......... .......... .......... 66%  102M 1s
 15450K .......... .......... .......... .......... .......... 67%  138M 1s
 15500K .......... .......... .......... .......... .......... 67% 71.8M 1s
 15550K .......... .......... .......... .......... .......... 67% 25.9M 1s
 15600K .......... .......... .......... .......... .......... 67%  108M 1s
 15650K .......... .......... .......... .......... .......... 68%  110M 1s
 15700K .......... .......... .......... .......... .......... 68%  138M 1s
 15750K .......... .......... .......... .......... .......... 68% 84.4M 1s
 15800K .......... .......... .......... .......... .......... 68%  144M 1s
 15850K .......... .......... .......... .......... .......... 68%  115M 1s
 15900K .......... .......... .......... .......... .......... 69%  109M 1s
 15950K .......... .......... .......... .......... .......... 69%  108M 1s
 16000K .......... .......... .......... .......... .......... 69%  173M 1s
 16050K .......... .......... .......... .......... .......... 69%  143M 1s
 16100K .......... .......... .......... .......... .......... 70% 98.0M 1s
 16150K .......... .......... .......... .......... .......... 70%  140M 1s
 16200K .......... .......... .......... .......... .......... 70% 99.9M 1s
 16250K .......... .......... .......... .......... .......... 70%  165M 1s
 16300K .......... .......... .......... .......... .......... 70% 95.4M 1s
 16350K .......... .......... .......... .......... .......... 71%  103M 1s
 16400K .......... .......... .......... .......... .......... 71% 97.7M 1s
 16450K .......... .......... .......... .......... .......... 71%  431M 1s
 16500K .......... .......... .......... .......... .......... 71% 96.6M 1s
 16550K .......... .......... .......... .......... .......... 71%  104M 1s
 16600K .......... .......... .......... .......... .......... 72%  199M 1s
 16650K .......... .......... .......... .......... .......... 72% 90.0M 1s
 16700K .......... .......... .......... .......... .......... 72%  124M 1s
 16750K .......... .......... .......... .......... .......... 72%  177M 1s
 16800K .......... .......... .......... .......... .......... 73% 81.4M 1s
 16850K .......... .......... .......... .......... .......... 73%  838M 1s
 16900K .......... .......... .......... .......... .......... 73% 85.5M 1s
 16950K .......... .......... .......... .......... .......... 73%  108M 1s
 17000K .......... .......... .......... .......... .......... 73% 74.2M 1s
 17050K .......... .......... .......... .......... .......... 74% 27.3M 1s
 17100K .......... .......... .......... .......... .......... 74%  437M 1s
 17150K .......... .......... .......... .......... .......... 74%  724M 1s
 17200K .......... .......... .......... .......... .......... 74% 67.0M 1s
 17250K .......... .......... .......... .......... .......... 74% 76.8M 1s
 17300K .......... .......... .......... .......... .......... 75% 79.4M 1s
 17350K .......... .......... .......... .......... .......... 75% 63.5M 1s
 17400K .......... .......... .......... .......... .......... 75% 62.6M 1s
 17450K .......... .......... .......... .......... .......... 75%  106M 1s
 17500K .......... .......... .......... .......... .......... 76% 71.3M 1s
 17550K .......... .......... .......... .......... .......... 76% 72.7M 1s
 17600K .......... .......... .......... .......... .......... 76% 79.7M 1s
 17650K .......... .......... .......... .......... .......... 76% 61.3M 1s
 17700K .......... .......... .......... .......... .......... 76% 83.8M 1s
 17750K .......... .......... .......... .......... .......... 77% 57.2M 1s
 17800K .......... .......... .......... .......... .......... 77% 72.8M 1s
 17850K .......... .......... .......... .......... .......... 77% 85.3M 1s
 17900K .......... .......... .......... .......... .......... 77% 75.9M 1s
 17950K .......... .......... .......... .......... .......... 78% 79.9M 1s
 18000K .......... .......... .......... .......... .......... 78% 74.7M 1s
 18050K .......... .......... .......... .......... .......... 78% 72.3M 1s
 18100K .......... .......... .......... .......... .......... 78% 71.6M 1s
 18150K .......... .......... .......... .......... .......... 78% 74.1M 1s
 18200K .......... .......... .......... .......... .......... 79% 70.8M 1s
 18250K .......... .......... .......... .......... .......... 79% 58.5M 1s
 18300K .......... .......... .......... .......... .......... 79% 30.2M 1s
 18350K .......... .......... .......... .......... .......... 79% 2.97G 1s
 18400K .......... .......... .......... .......... .......... 79%  272M 0s
 18450K .......... .......... .......... .......... .......... 80% 70.0M 0s
 18500K .......... .......... .......... .......... .......... 80% 74.9M 0s
 18550K .......... .......... .......... .......... .......... 80% 75.4M 0s
 18600K .......... .......... .......... .......... .......... 80% 60.4M 0s
 18650K .......... .......... .......... .......... .......... 81% 88.7M 0s
 18700K .......... .......... .......... .......... .......... 81% 76.0M 0s
 18750K .......... .......... .......... .......... .......... 81% 71.4M 0s
 18800K .......... .......... .......... .......... .......... 81% 65.9M 0s
 18850K .......... .......... .......... .......... .......... 81% 68.7M 0s
 18900K .......... .......... .......... .......... .......... 82% 67.3M 0s
 18950K .......... .......... .......... .......... .......... 82% 29.0M 0s
 19000K .......... .......... .......... .......... .......... 82% 94.1M 0s
 19050K .......... .......... .......... .......... .......... 82%  109M 0s
 19100K .......... .......... .......... .......... .......... 83% 74.7M 0s
 19150K .......... .......... .......... .......... .......... 83%  131M 0s
 19200K .......... .......... .......... .......... .......... 83% 58.5M 0s
 19250K .......... .......... .......... .......... .......... 83% 83.3M 0s
 19300K .......... .......... .......... .......... .......... 83%  103M 0s
 19350K .......... .......... .......... .......... .......... 84%  108M 0s
 19400K .......... .......... .......... .......... .......... 84%  104M 0s
 19450K .......... .......... .......... .......... .......... 84% 69.2M 0s
 19500K .......... .......... .......... .......... .......... 84% 71.1M 0s
 19550K .......... .......... .......... .......... .......... 84% 77.0M 0s
 19600K .......... .......... .......... .......... .......... 85% 79.4M 0s
 19650K .......... .......... .......... .......... .......... 85% 66.7M 0s
 19700K .......... .......... .......... .......... .......... 85% 73.1M 0s
 19750K .......... .......... .......... .......... .......... 85% 52.9M 0s
 19800K .......... .......... .......... .......... .......... 86% 10.9M 0s
 19850K .......... .......... .......... .......... .......... 86% 82.0M 0s
 19900K .......... .......... .......... .......... .......... 86% 82.5M 0s
 19950K .......... .......... .......... .......... .......... 86%  113M 0s
 20000K .......... .......... .......... .......... .......... 86%  114M 0s
 20050K .......... .......... .......... .......... .......... 87% 94.7M 0s
 20100K .......... .......... .......... .......... .......... 87% 21.7M 0s
 20150K .......... .......... .......... .......... .......... 87%  290M 0s
 20200K .......... .......... .......... .......... .......... 87% 83.4M 0s
 20250K .......... .......... .......... .......... .......... 87% 93.7M 0s
 20300K .......... .......... .......... .......... .......... 88%  121M 0s
 20350K .......... .......... .......... .......... .......... 88%  118M 0s
 20400K .......... .......... .......... .......... .......... 88%  122M 0s
 20450K .......... .......... .......... .......... .......... 88%  135M 0s
 20500K .......... .......... .......... .......... .......... 89%  122M 0s
 20550K .......... .......... .......... .......... .......... 89%  114M 0s
 20600K .......... .......... .......... .......... .......... 89%  102M 0s
 20650K .......... .......... .......... .......... .......... 89% 97.9M 0s
 20700K .......... .......... .......... .......... .......... 89%  154M 0s
 20750K .......... .......... .......... .......... .......... 90% 90.9M 0s
 20800K .......... .......... .......... .......... .......... 90%  247M 0s
 20850K .......... .......... .......... .......... .......... 90% 93.2M 0s
 20900K .......... .......... .......... .......... .......... 90% 91.9M 0s
 20950K .......... .......... .......... .......... .......... 91% 95.3M 0s
 21000K .......... .......... .......... .......... .......... 91%  210M 0s
 21050K .......... .......... .......... .......... .......... 91% 85.1M 0s
 21100K .......... .......... .......... .......... .......... 91%  103M 0s
 21150K .......... .......... .......... .......... .......... 91% 84.3M 0s
 21200K .......... .......... .......... .......... .......... 92% 29.3M 0s
 21250K .......... .......... .......... .......... .......... 92% 2.11G 0s
 21300K .......... .......... .......... .......... .......... 92%  111M 0s
 21350K .......... .......... .......... .......... .......... 92% 81.9M 0s
 21400K .......... .......... .......... .......... .......... 92% 79.8M 0s
 21450K .......... .......... .......... .......... .......... 93% 64.9M 0s
 21500K .......... .......... .......... .......... .......... 93% 79.9M 0s
 21550K .......... .......... .......... .......... .......... 93% 70.4M 0s
 21600K .......... .......... .......... .......... .......... 93% 57.1M 0s
 21650K .......... .......... .......... .......... .......... 94% 97.7M 0s
 21700K .......... .......... .......... .......... .......... 94% 86.5M 0s
 21750K .......... .......... .......... .......... .......... 94% 57.6M 0s
 21800K .......... .......... .......... .......... .......... 94% 70.5M 0s
 21850K .......... .......... .......... .......... .......... 94% 78.7M 0s
 21900K .......... .......... .......... .......... .......... 95% 91.0M 0s
 21950K .......... .......... .......... .......... .......... 95% 72.4M 0s
 22000K .......... .......... .......... .......... .......... 95% 63.0M 0s
 22050K .......... .......... .......... .......... .......... 95% 71.0M 0s
 22100K .......... .......... .......... .......... .......... 96% 88.1M 0s
 22150K .......... .......... .......... .......... .......... 96% 73.3M 0s
 22200K .......... .......... .......... .......... .......... 96% 77.1M 0s
 22250K .......... .......... .......... .......... .......... 96% 74.8M 0s
 22300K .......... .......... .......... .......... .......... 96% 72.9M 0s
 22350K .......... .......... .......... .......... .......... 97% 63.1M 0s
 22400K .......... .......... .......... .......... .......... 97% 77.3M 0s
 22450K .......... .......... .......... .......... .......... 97% 13.5M 0s
 22500K .......... .......... .......... .......... .......... 97% 48.3M 0s
 22550K .......... .......... .......... .......... .......... 97% 41.3M 0s
 22600K .......... .......... .......... .......... .......... 98% 55.9M 0s
 22650K .......... .......... .......... .......... .......... 98% 68.4M 0s
 22700K .......... .......... .......... .......... .......... 98% 59.7M 0s
 22750K .......... .......... .......... .......... .......... 98% 83.9M 0s
 22800K .......... .......... .......... .......... .......... 99% 70.4M 0s
 22850K .......... .......... .......... .......... .......... 99% 69.2M 0s
 22900K .......... .......... .......... .......... .......... 99% 96.8M 0s
 22950K .......... .......... .......... .......... .......... 99%  108M 0s
 23000K .......... .......... .......... .......... .......... 99% 73.0M 0s
 23050K .......... ........                                   100% 96.1M=2.5s

2020-03-02 03:24:16 (74.7 Mb/s) - ‘/dev/null’ saved [23622382/23622382]

