--2020-02-25 22:14:14--  http://www.comures.org.sv/CIRCULAR-043-2017.pdf%0D
Resolving www.comures.org.sv (www.comures.org.sv)... 174.142.89.94
Connecting to www.comures.org.sv (www.comures.org.sv)|174.142.89.94|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:15 ERROR 404: Not Found.

--2020-02-25 22:14:39--  http://www.comures.org.sv/CIRCULAR-043-2017.pdf%0D
Resolving www.comures.org.sv (www.comures.org.sv)... 174.142.89.94
Connecting to www.comures.org.sv (www.comures.org.sv)|174.142.89.94|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:39 ERROR 404: Not Found.

