--2020-02-25 22:13:53--  http://biblioteca.utec.edu.sv/siab/virtual/DiarioOficial/publicaciones2004/enero/20040116S.pdf%0D
Resolving biblioteca.utec.edu.sv (biblioteca.utec.edu.sv)... 181.225.132.82
Connecting to biblioteca.utec.edu.sv (biblioteca.utec.edu.sv)|181.225.132.82|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:54 ERROR 404: Not Found.

--2020-02-25 22:14:20--  http://biblioteca.utec.edu.sv/siab/virtual/DiarioOficial/publicaciones2004/enero/20040116S.pdf%0D
Resolving biblioteca.utec.edu.sv (biblioteca.utec.edu.sv)... 181.225.132.82
Connecting to biblioteca.utec.edu.sv (biblioteca.utec.edu.sv)|181.225.132.82|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:20 ERROR 404: Not Found.

