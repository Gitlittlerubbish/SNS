--2020-02-25 22:12:51--  https://www.tsc.gob.sv/pdf/constitucionsv.pdf%0D
Resolving www.tsc.gob.sv (www.tsc.gob.sv)... 104.27.170.247, 104.27.171.247
Connecting to www.tsc.gob.sv (www.tsc.gob.sv)|104.27.170.247|:443... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:12:52 ERROR 404: Not Found.

--2020-02-25 22:13:28--  https://www.tsc.gob.sv/pdf/constitucionsv.pdf%0D
Resolving www.tsc.gob.sv (www.tsc.gob.sv)... 104.27.171.247, 104.27.170.247
Connecting to www.tsc.gob.sv (www.tsc.gob.sv)|104.27.171.247|:443... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:28 ERROR 404: Not Found.

