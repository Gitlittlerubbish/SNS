--2020-02-25 22:12:43--  https://www.transparencia.gob.sv/institutions/isss/documents/7853/download%0D
Resolving www.transparencia.gob.sv (www.transparencia.gob.sv)... 95.216.118.177
Connecting to www.transparencia.gob.sv (www.transparencia.gob.sv)|95.216.118.177|:443... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:12:43 ERROR 404: Not Found.

--2020-02-25 22:13:22--  https://www.transparencia.gob.sv/institutions/isss/documents/7853/download%0D
Resolving www.transparencia.gob.sv (www.transparencia.gob.sv)... 95.216.118.177
Connecting to www.transparencia.gob.sv (www.transparencia.gob.sv)|95.216.118.177|:443... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:23 ERROR 404: Not Found.

