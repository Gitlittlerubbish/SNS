--2020-03-02 03:27:26--  http://www.censos.gob.sv/cpv/descargas/CPV_Proyeccion_Resultados.pdf
Resolving www.censos.gob.sv (www.censos.gob.sv)... 200.89.85.145
Connecting to www.censos.gob.sv (www.censos.gob.sv)|200.89.85.145|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 446731 (436K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 11%  676K 5s
    50K .......... .......... .......... .......... .......... 22% 2.66M 3s
   100K .......... .......... .......... .......... .......... 34% 32.7M 1s
   150K .......... .......... .......... .......... .......... 45% 2.90M 1s
   200K .......... .......... .......... .......... .......... 57%  102M 1s
   250K .......... .......... .......... .......... .......... 68% 4.23M 0s
   300K .......... .......... .......... .......... .......... 80% 7.58M 0s
   350K .......... .......... .......... .......... .......... 91%  141M 0s
   400K .......... .......... .......... ......               100%  106M=1.1s

2020-03-02 03:27:27 (3.33 Mb/s) - ‘/dev/null’ saved [446731/446731]

