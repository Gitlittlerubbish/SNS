--2020-03-02 03:25:57--  http://ovisss.isss.gob.sv/documentos_ofivi/Calendario_OVISSS_2020.pdf
Resolving ovisss.isss.gob.sv (ovisss.isss.gob.sv)... 129.158.125.97
Connecting to ovisss.isss.gob.sv (ovisss.isss.gob.sv)|129.158.125.97|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: https://ovisss.isss.gob.sv/documentos_ofivi/Calendario_OVISSS_2020.pdf [following]
--2020-03-02 03:25:58--  https://ovisss.isss.gob.sv/documentos_ofivi/Calendario_OVISSS_2020.pdf
Connecting to ovisss.isss.gob.sv (ovisss.isss.gob.sv)|129.158.125.97|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: 420045 (410K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 12%  695K 4s
    50K .......... .......... .......... .......... .......... 24%  571K 4s
   100K .......... .......... .......... .......... .......... 36%  330M 2s
   150K .......... .......... .......... .......... .......... 48%  278K 3s
   200K .......... .......... .......... .......... .......... 60%  664M 2s
   250K .......... .......... .......... .......... .......... 73%  520K 1s
   300K .......... .......... .......... .......... .......... 85% 10.3M 1s
   350K .......... .......... .......... .......... .......... 97%  470K 0s
   400K ..........                                            100% 1.61G=4.5s

2020-03-02 03:26:05 (750 Kb/s) - ‘/dev/null’ saved [420045/420045]

