--2020-03-02 03:23:41--  http://www.transparenciafiscal.gob.sv/downloads/pdf/DC5544_CAP_21.pdf
Resolving www.transparenciafiscal.gob.sv (www.transparenciafiscal.gob.sv)... 190.5.131.23, 190.57.24.31
Connecting to www.transparenciafiscal.gob.sv (www.transparenciafiscal.gob.sv)|190.5.131.23|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 19989 (20K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .........                                  100%  560K=0.3s

2020-03-02 03:23:42 (560 Kb/s) - ‘/dev/null’ saved [19989/19989]

