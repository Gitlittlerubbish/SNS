--2020-03-02 03:25:52--  http://www.minsal.sv/archivos/chagas2008/pdf/La_enfermedad_de_chagas_en_el_salvador_evolucion_historica_y_desafio_para_el_control.pdf
Resolving www.minsal.sv (www.minsal.sv)... 190.86.223.123
Connecting to www.minsal.sv (www.minsal.sv)|190.86.223.123|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 4491613 (4.3M) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  1% 1.52M 23s
    50K .......... .......... .......... .......... ..........  2% 2.96M 17s
   100K .......... .......... .......... .......... ..........  3%  228M 12s
   150K .......... .......... .......... .......... ..........  4% 96.1M 9s
   200K .......... .......... .......... .......... ..........  5% 2.62M 9s
   250K .......... .......... .......... .......... ..........  6%  124M 8s
   300K .......... .......... .......... .......... ..........  7% 3.74M 8s
   350K .......... .......... .......... .......... ..........  9%  104M 7s
   400K .......... .......... .......... .......... .......... 10% 2.98M 7s
   450K .......... .......... .......... .......... .......... 11% 1.42G 6s
   500K .......... .......... .......... .......... .......... 12% 1.27G 6s
   550K .......... .......... .......... .......... .......... 13% 1.53G 5s
   600K .......... .......... .......... .......... .......... 14% 1.53G 5s
   650K .......... .......... .......... .......... .......... 15% 3.02M 5s
   700K .......... .......... .......... .......... .......... 17% 2.92M 5s
   750K .......... .......... .......... .......... .......... 18% 1.36G 5s
   800K .......... .......... .......... .......... .......... 19%  108M 5s
   850K .......... .......... .......... .......... .......... 20% 2.06G 4s
   900K .......... .......... .......... .......... .......... 21% 1.65G 4s
   950K .......... .......... .......... .......... .......... 22% 3.16M 4s
  1000K .......... .......... .......... .......... .......... 23%  123M 4s
  1050K .......... .......... .......... .......... .......... 25% 2.95M 4s
  1100K .......... .......... .......... .......... .......... 26% 1.43G 4s
  1150K .......... .......... .......... .......... .......... 27%  431M 4s
  1200K .......... .......... .......... .......... .......... 28% 1.23G 3s
  1250K .......... .......... .......... .......... .......... 29% 3.09M 4s
  1300K .......... .......... .......... .......... .......... 30%  243M 3s
  1350K .......... .......... .......... .......... .......... 31%  234M 3s
  1400K .......... .......... .......... .......... .......... 33% 3.06M 3s
  1450K .......... .......... .......... .......... .......... 34%  206M 3s
  1500K .......... .......... .......... .......... .......... 35%  203M 3s
  1550K .......... .......... .......... .......... .......... 36% 3.10M 3s
  1600K .......... .......... .......... .......... .......... 37%  144M 3s
  1650K .......... .......... .......... .......... .......... 38%  120M 3s
  1700K .......... .......... .......... .......... .......... 39% 3.19M 3s
  1750K .......... .......... .......... .......... .......... 41%  141M 3s
  1800K .......... .......... .......... .......... .......... 42%  117M 3s
  1850K .......... .......... .......... .......... .......... 43% 3.18M 3s
  1900K .......... .......... .......... .......... .......... 44%  104M 3s
  1950K .......... .......... .......... .......... .......... 45% 92.9M 2s
  2000K .......... .......... .......... .......... .......... 46%  463M 2s
  2050K .......... .......... .......... .......... .......... 47% 3.16M 2s
  2100K .......... .......... .......... .......... .......... 49% 91.6M 2s
  2150K .......... .......... .......... .......... .......... 50%  204M 2s
  2200K .......... .......... .......... .......... .......... 51% 3.17M 2s
  2250K .......... .......... .......... .......... .......... 52% 96.7M 2s
  2300K .......... .......... .......... .......... .......... 53%  114M 2s
  2350K .......... .......... .......... .......... .......... 54% 3.31M 2s
  2400K .......... .......... .......... .......... .......... 55% 92.6M 2s
  2450K .......... .......... .......... .......... .......... 56%  108M 2s
  2500K .......... .......... .......... .......... .......... 58% 3.36M 2s
  2550K .......... .......... .......... .......... .......... 59% 38.2M 2s
  2600K .......... .......... .......... .......... .......... 60%  130M 2s
  2650K .......... .......... .......... .......... .......... 61% 3.49M 2s
  2700K .......... .......... .......... .......... .......... 62% 27.3M 2s
  2750K .......... .......... .......... .......... .......... 63%  222M 2s
  2800K .......... .......... .......... .......... .......... 64%  111M 1s
  2850K .......... .......... .......... .......... .......... 66% 3.18M 1s
  2900K .......... .......... .......... .......... .......... 67%  163M 1s
  2950K .......... .......... .......... .......... .......... 68%  148M 1s
  3000K .......... .......... .......... .......... .......... 69% 3.41M 1s
  3050K .......... .......... .......... .......... .......... 70% 29.3M 1s
  3100K .......... .......... .......... .......... .......... 71%  356M 1s
  3150K .......... .......... .......... .......... .......... 72% 3.55M 1s
  3200K .......... .......... .......... .......... .......... 74% 22.8M 1s
  3250K .......... .......... .......... .......... .......... 75%  119M 1s
  3300K .......... .......... .......... .......... .......... 76%  232M 1s
  3350K .......... .......... .......... .......... .......... 77% 1.56M 1s
  3400K .......... .......... .......... .......... .......... 78% 1.65G 1s
  3450K .......... .......... .......... .......... .......... 79% 1.69G 1s
  3500K .......... .......... .......... .......... .......... 80% 1.99G 1s
  3550K .......... .......... .......... .......... .......... 82%  111M 1s
  3600K .......... .......... .......... .......... .......... 83% 3.60M 1s
  3650K .......... .......... .......... .......... .......... 84% 22.6M 1s
  3700K .......... .......... .......... .......... .......... 85% 84.6M 1s
  3750K .......... .......... .......... .......... .......... 86% 3.38M 1s
  3800K .......... .......... .......... .......... .......... 87% 37.3M 1s
  3850K .......... .......... .......... .......... .......... 88% 3.62M 0s
  3900K .......... .......... .......... .......... .......... 90% 22.6M 0s
  3950K .......... .......... .......... .......... .......... 91% 73.3M 0s
  4000K .......... .......... .......... .......... .......... 92% 3.44M 0s
  4050K .......... .......... .......... .......... .......... 93% 34.7M 0s
  4100K .......... .......... .......... .......... .......... 94% 80.5M 0s
  4150K .......... .......... .......... .......... .......... 95% 3.38M 0s
  4200K .......... .......... .......... .......... .......... 96% 41.0M 0s
  4250K .......... .......... .......... .......... .......... 98% 3.63M 0s
  4300K .......... .......... .......... .......... .......... 99% 25.6M 0s
  4350K .......... .......... .......... ......               100% 56.9M=4.2s

2020-03-02 03:25:57 (8.51 Mb/s) - ‘/dev/null’ saved [4491613/4491613]

