--2020-02-25 22:14:01--  https://www.bolsadevalores.com.sv/files/29027/FF_OPTIMASERVICIOSFINANCIEROS_201812_PCR.pdf%0D
Resolving www.bolsadevalores.com.sv (www.bolsadevalores.com.sv)... 190.5.141.232
Connecting to www.bolsadevalores.com.sv (www.bolsadevalores.com.sv)|190.5.141.232|:443... connected.
HTTP request sent, awaiting response... 403 Forbidden
2020-02-25 22:14:02 ERROR 403: Forbidden.

--2020-02-25 22:14:28--  https://www.bolsadevalores.com.sv/files/29027/FF_OPTIMASERVICIOSFINANCIEROS_201812_PCR.pdf%0D
Resolving www.bolsadevalores.com.sv (www.bolsadevalores.com.sv)... 190.5.141.232
Connecting to www.bolsadevalores.com.sv (www.bolsadevalores.com.sv)|190.5.141.232|:443... connected.
HTTP request sent, awaiting response... 403 Forbidden
2020-02-25 22:14:28 ERROR 403: Forbidden.

