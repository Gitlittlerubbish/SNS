--2020-02-25 22:12:48--  https://unasa.edu.sv/PDF/cat%25C3%25A1logo_2018_UNASA.pdf%0D
Resolving unasa.edu.sv (unasa.edu.sv)... 74.220.199.65
Connecting to unasa.edu.sv (unasa.edu.sv)|74.220.199.65|:443... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:12:49 ERROR 404: Not Found.

--2020-02-25 22:13:25--  https://unasa.edu.sv/PDF/cat%25C3%25A1logo_2018_UNASA.pdf%0D
Resolving unasa.edu.sv (unasa.edu.sv)... 74.220.199.65
Connecting to unasa.edu.sv (unasa.edu.sv)|74.220.199.65|:443... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:26 ERROR 404: Not Found.

