--2020-02-25 22:13:39--  http://aplicaciones.itca.edu.sv/PwdCorreoITCA.pdf%0D
Resolving aplicaciones.itca.edu.sv (aplicaciones.itca.edu.sv)... 200.35.188.115
Connecting to aplicaciones.itca.edu.sv (aplicaciones.itca.edu.sv)|200.35.188.115|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:40 ERROR 404: Not Found.

--2020-02-25 22:14:09--  http://aplicaciones.itca.edu.sv/PwdCorreoITCA.pdf%0D
Resolving aplicaciones.itca.edu.sv (aplicaciones.itca.edu.sv)... 200.35.188.115
Connecting to aplicaciones.itca.edu.sv (aplicaciones.itca.edu.sv)|200.35.188.115|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:14:10 ERROR 404: Not Found.

