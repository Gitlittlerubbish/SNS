--2020-02-25 22:12:53--  http://www.jurisprudencia.gob.sv/publicados/Juris_Publicados_Junio2019v3.pdf%0D
Resolving www.jurisprudencia.gob.sv (www.jurisprudencia.gob.sv)... 200.31.169.67
Connecting to www.jurisprudencia.gob.sv (www.jurisprudencia.gob.sv)|200.31.169.67|:80... connected.
HTTP request sent, awaiting response... 403 Forbidden
2020-02-25 22:12:53 ERROR 403: Forbidden.

--2020-02-25 22:13:29--  http://www.jurisprudencia.gob.sv/publicados/Juris_Publicados_Junio2019v3.pdf%0D
Resolving www.jurisprudencia.gob.sv (www.jurisprudencia.gob.sv)... 200.31.169.67
Connecting to www.jurisprudencia.gob.sv (www.jurisprudencia.gob.sv)|200.31.169.67|:80... connected.
HTTP request sent, awaiting response... 403 Forbidden
2020-02-25 22:13:29 ERROR 403: Forbidden.

