--2020-02-25 22:12:54--  http://www.amate.org.sv/doc/LGBT_Shadow_Report_El_Salvador_HRC100.pdf%0D
Resolving www.amate.org.sv (www.amate.org.sv)... 107.180.51.78
Connecting to www.amate.org.sv (www.amate.org.sv)|107.180.51.78|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K .......... .......... ....                             1.62M=0.1s

2020-02-25 22:12:54 (1.62 Mb/s) - ‘/dev/null’ saved [24850]

--2020-02-25 22:12:54--  http://www.amate.org.sv/doc/LGBT_Shadow_Report_El_Salvador_HRC100.pdf%0D
Resolving www.amate.org.sv (www.amate.org.sv)... 107.180.51.78
Connecting to www.amate.org.sv (www.amate.org.sv)|107.180.51.78|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K .......... .......... ....                             1.63M=0.1s

2020-02-25 22:12:55 (1.63 Mb/s) - ‘/dev/null’ saved [24850]

--2020-02-25 22:13:30--  http://www.amate.org.sv/doc/LGBT_Shadow_Report_El_Salvador_HRC100.pdf%0D
Resolving www.amate.org.sv (www.amate.org.sv)... 107.180.51.78
Connecting to www.amate.org.sv (www.amate.org.sv)|107.180.51.78|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K .......... .......... ....                             2.25M=0.09s

2020-02-25 22:13:30 (2.25 Mb/s) - ‘/dev/null’ saved [24850]

--2020-02-25 22:13:30--  http://www.amate.org.sv/doc/LGBT_Shadow_Report_El_Salvador_HRC100.pdf%0D
Resolving www.amate.org.sv (www.amate.org.sv)... 107.180.51.78
Connecting to www.amate.org.sv (www.amate.org.sv)|107.180.51.78|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K .......... .......... ....                             1.96M=0.1s

2020-02-25 22:13:30 (1.96 Mb/s) - ‘/dev/null’ saved [24850]

