--2020-02-25 22:14:02--  https://tienda.movistar.com.sv/tv/Movistar_TvHD_Manual_Uso.pdf%0D
Resolving tienda.movistar.com.sv (tienda.movistar.com.sv)... 72.47.233.224
Connecting to tienda.movistar.com.sv (tienda.movistar.com.sv)|72.47.233.224|:443... connected.
HTTP request sent, awaiting response... 302 Found
Location: https://tienda.movistar.com.sv/404/ [following]
--2020-02-25 22:14:03--  https://tienda.movistar.com.sv/404/
Reusing existing connection to tienda.movistar.com.sv:443.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K ......                                                 2.19G=0s

2020-02-25 22:14:04 (2.19 Gb/s) - ‘/dev/null’ saved [6461]

--2020-02-25 22:14:04--  https://tienda.movistar.com.sv/tv/Movistar_TvHD_Manual_Uso.pdf%0D
Resolving tienda.movistar.com.sv (tienda.movistar.com.sv)... 72.47.233.224
Connecting to tienda.movistar.com.sv (tienda.movistar.com.sv)|72.47.233.224|:443... connected.
HTTP request sent, awaiting response... 302 Found
Location: https://tienda.movistar.com.sv/404/ [following]
--2020-02-25 22:14:04--  https://tienda.movistar.com.sv/404/
Reusing existing connection to tienda.movistar.com.sv:443.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K ......                                                 1.78G=0s

2020-02-25 22:14:04 (1.78 Gb/s) - ‘/dev/null’ saved [6461]

--2020-02-25 22:14:28--  https://tienda.movistar.com.sv/tv/Movistar_TvHD_Manual_Uso.pdf%0D
Resolving tienda.movistar.com.sv (tienda.movistar.com.sv)... 72.47.233.224
Connecting to tienda.movistar.com.sv (tienda.movistar.com.sv)|72.47.233.224|:443... connected.
HTTP request sent, awaiting response... 302 Found
Location: https://tienda.movistar.com.sv/404/ [following]
--2020-02-25 22:14:29--  https://tienda.movistar.com.sv/404/
Reusing existing connection to tienda.movistar.com.sv:443.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K ......                                                 1.03G=0s

2020-02-25 22:14:29 (1.03 Gb/s) - ‘/dev/null’ saved [6461]

--2020-02-25 22:14:29--  https://tienda.movistar.com.sv/tv/Movistar_TvHD_Manual_Uso.pdf%0D
Resolving tienda.movistar.com.sv (tienda.movistar.com.sv)... 72.47.233.224
Connecting to tienda.movistar.com.sv (tienda.movistar.com.sv)|72.47.233.224|:443... connected.
HTTP request sent, awaiting response... 302 Found
Location: https://tienda.movistar.com.sv/404/ [following]
--2020-02-25 22:14:30--  https://tienda.movistar.com.sv/404/
Reusing existing connection to tienda.movistar.com.sv:443.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K ......                                                 2.23G=0s

2020-02-25 22:14:30 (2.23 Gb/s) - ‘/dev/null’ saved [6461]

