--2020-03-02 03:23:36--  http://biblioteca.ues.edu.sv/revistas/10800099.pdf
Resolving biblioteca.ues.edu.sv (biblioteca.ues.edu.sv)... 168.232.48.132
Connecting to biblioteca.ues.edu.sv (biblioteca.ues.edu.sv)|168.232.48.132|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 320589 (313K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 15%  651K 3s
    50K .......... .......... .......... .......... .......... 31% 1.30M 2s
   100K .......... .......... .......... .......... .......... 47% 2.61M 1s
   150K .......... .......... .......... .......... .......... 63%  130M 1s
   200K .......... .......... .......... .......... .......... 79% 2.62M 0s
   250K .......... .......... .......... .......... .......... 95% 4.20M 0s
   300K .......... ...                                        100% 1.84M=1.4s

2020-03-02 03:23:39 (1.81 Mb/s) - ‘/dev/null’ saved [320589/320589]

--2020-03-02 03:23:39--  http://biblioteca.ues.edu.sv/revistas/10800057E1.pdf
Resolving biblioteca.ues.edu.sv (biblioteca.ues.edu.sv)... 168.232.48.132
Connecting to biblioteca.ues.edu.sv (biblioteca.ues.edu.sv)|168.232.48.132|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 370301 (362K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 13%  653K 4s
    50K .......... .......... .......... .......... .......... 27% 2.59M 2s
   100K .......... .......... .......... .......... .......... 41% 2.58M 1s
   150K .......... .......... .......... .......... .......... 55% 2.60M 1s
   200K .......... .......... .......... .......... .......... 69% 2.63M 1s
   250K .......... .......... .......... .......... .......... 82%  155M 0s
   300K .......... .......... .......... .......... .......... 96% 2.70M 0s
   350K .......... .                                          100%  105M=1.4s

2020-03-02 03:23:41 (2.10 Mb/s) - ‘/dev/null’ saved [370301/370301]

