--2020-02-25 22:12:52--  https://www.fomilenioii.gob.sv/asset/documents/90%0D
Resolving www.fomilenioii.gob.sv (www.fomilenioii.gob.sv)... 138.201.55.180
Connecting to www.fomilenioii.gob.sv (www.fomilenioii.gob.sv)|138.201.55.180|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [application/x-download]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 6.81M
    50K .......... .......... .......... .......... .......... 16.8M
   100K .......... .......... .......... .......... .......... 1.33G
   150K .......... .......... .......... .......... .......... 17.0M
   200K .......... .......... .......... .......... ..........  405M
   250K .......... .......... .......... .......... ..........  386M
   300K .......... .......... .......... .......... .......... 1.99G
   350K .......... .......... .......... .......... .......... 18.3M
   400K .......... .......... .......... .......... .......... 1.03G
   450K .......... .......... .                                 421M=0.1s

2020-02-25 22:12:53 (28.8 Mb/s) - ‘/dev/null’ saved [482980]

--2020-02-25 22:12:53--  https://www.fomilenioii.gob.sv/asset/documents/90%0D
Resolving www.fomilenioii.gob.sv (www.fomilenioii.gob.sv)... 138.201.55.180
Connecting to www.fomilenioii.gob.sv (www.fomilenioii.gob.sv)|138.201.55.180|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [application/x-download]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 8.30M
    50K .......... .......... .......... .......... .......... 17.3M
   100K .......... .......... .......... .......... ..........  518M
   150K .......... .......... .......... .......... .......... 17.3M
   200K .......... .......... .......... .......... ..........  698M
   250K .......... .......... .......... .......... ..........  829M
   300K .......... .......... .......... .......... ..........  768M
   350K .......... .......... .......... .......... .......... 17.4M
   400K .......... .......... .......... .......... ..........  449M
   450K .......... .......... .                                 786M=0.1s

2020-02-25 22:12:53 (31.2 Mb/s) - ‘/dev/null’ saved [482980]

--2020-02-25 22:13:28--  https://www.fomilenioii.gob.sv/asset/documents/90%0D
Resolving www.fomilenioii.gob.sv (www.fomilenioii.gob.sv)... 138.201.55.180
Connecting to www.fomilenioii.gob.sv (www.fomilenioii.gob.sv)|138.201.55.180|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [application/x-download]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 8.42M
    50K .......... .......... .......... .......... .......... 16.7M
   100K .......... .......... .......... .......... ..........  112M
   150K .......... .......... .......... .......... .......... 19.5M
   200K .......... .......... .......... .......... ..........  394M
   250K .......... .......... .......... .......... ..........  139M
   300K .......... .......... .......... .......... .......... 20.9M
   350K .......... .......... .......... .......... ..........  564M
   400K .......... .......... .......... .......... ..........  369M
   450K .......... .......... .                                 455M=0.1s

2020-02-25 22:13:29 (31.3 Mb/s) - ‘/dev/null’ saved [482980]

--2020-02-25 22:13:29--  https://www.fomilenioii.gob.sv/asset/documents/90%0D
Resolving www.fomilenioii.gob.sv (www.fomilenioii.gob.sv)... 138.201.55.180
Connecting to www.fomilenioii.gob.sv (www.fomilenioii.gob.sv)|138.201.55.180|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [application/x-download]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 8.34M
    50K .......... .......... .......... .......... .......... 16.5M
   100K .......... .......... .......... .......... .......... 3.42G
   150K .......... .......... .......... .......... .......... 17.0M
   200K .......... .......... .......... .......... ..........  358M
   250K .......... .......... .......... .......... ..........  403M
   300K .......... .......... .......... .......... .......... 18.7M
   350K .......... .......... .......... .......... .......... 2.73G
   400K .......... .......... .......... .......... ..........  603M
   450K .......... .......... .                                 406M=0.1s

2020-02-25 22:13:29 (31.3 Mb/s) - ‘/dev/null’ saved [482980]

