--2020-03-02 03:24:06--  http://www.integral.com.sv/asset/documents/859
Resolving www.integral.com.sv (www.integral.com.sv)... 95.216.241.9
Connecting to www.integral.com.sv (www.integral.com.sv)|95.216.241.9|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: https://www.integral.com.sv/asset/documents/859 [following]
--2020-03-02 03:24:06--  https://www.integral.com.sv/asset/documents/859
Connecting to www.integral.com.sv (www.integral.com.sv)|95.216.241.9|:443... connected.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 5.37M
    50K .......... .......... .......... ....                   315M=0.08s

2020-03-02 03:24:07 (8.94 Mb/s) - ‘/dev/null’ saved [86155]

