--2020-03-02 03:24:26--  http://www.amate.org.sv/doc/LGBT_Shadow_Report_El_Salvador_HRC100.pdf
Resolving www.amate.org.sv (www.amate.org.sv)... 107.180.51.78
Connecting to www.amate.org.sv (www.amate.org.sv)|107.180.51.78|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 344448 (336K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 14% 2.22M 1s
    50K .......... .......... .......... .......... .......... 29% 4.68M 1s
   100K .......... .......... .......... .......... .......... 44% 4.93M 0s
   150K .......... .......... .......... .......... .......... 59% 5.62M 0s
   200K .......... .......... .......... .......... .......... 74% 33.5M 0s
   250K .......... .......... .......... .......... .......... 89% 5.85M 0s
   300K .......... .......... .......... ......               100% 29.5M=0.5s

2020-03-02 03:24:27 (5.29 Mb/s) - ‘/dev/null’ saved [344448/344448]

