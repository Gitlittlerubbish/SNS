--2020-03-02 03:24:07--  http://www.fundar.org.sv/referencias/pipilpots.pdf
Resolving www.fundar.org.sv (www.fundar.org.sv)... 190.120.10.123
Connecting to www.fundar.org.sv (www.fundar.org.sv)|190.120.10.123|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 3385841 (3.2M) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... ..........  1% 1.45M 18s
    50K .......... .......... .......... .......... ..........  3% 2.97M 13s
   100K .......... .......... .......... .......... ..........  4% 3.01M 12s
   150K .......... .......... .......... .......... ..........  6% 3.03M 11s
   200K .......... .......... .......... .......... ..........  7% 3.02M 10s
   250K .......... .......... .......... .......... ..........  9% 3.03M 10s
   300K .......... .......... .......... .......... .......... 10% 3.07M 9s
   350K .......... .......... .......... .......... .......... 12% 3.05M 9s
   400K .......... .......... .......... .......... .......... 13% 3.10M 9s
   450K .......... .......... .......... .......... .......... 15% 3.12M 8s
   500K .......... .......... .......... .......... .......... 16% 3.17M 8s
   550K .......... .......... .......... .......... .......... 18% 32.2M 7s
   600K .......... .......... .......... .......... .......... 19% 3.12M 7s
   650K .......... .......... .......... .......... .......... 21% 3.13M 7s
   700K .......... .......... .......... .......... .......... 22% 3.39M 7s
   750K .......... .......... .......... .......... .......... 24% 19.4M 6s
   800K .......... .......... .......... .......... .......... 25% 3.07M 6s
   850K .......... .......... .......... .......... .......... 27% 3.34M 6s
   900K .......... .......... .......... .......... .......... 28% 26.5M 6s
   950K .......... .......... .......... .......... .......... 30% 3.21M 6s
  1000K .......... .......... .......... .......... .......... 31% 50.0M 5s
  1050K .......... .......... .......... .......... .......... 33% 3.04M 5s
  1100K .......... .......... .......... .......... .......... 34% 82.9M 5s
  1150K .......... .......... .......... .......... .......... 36% 3.13M 5s
  1200K .......... .......... .......... .......... .......... 37% 4.04M 5s
  1250K .......... .......... .......... .......... .......... 39% 12.4M 4s
  1300K .......... .......... .......... .......... .......... 40% 51.6M 4s
  1350K .......... .......... .......... .......... .......... 42% 3.26M 4s
  1400K .......... .......... .......... .......... .......... 43% 44.0M 4s
  1450K .......... .......... .......... .......... .......... 45% 3.32M 4s
  1500K .......... .......... .......... .......... .......... 46% 37.1M 4s
  1550K .......... .......... .......... .......... .......... 48% 3.36M 3s
  1600K .......... .......... .......... .......... .......... 49% 40.8M 3s
  1650K .......... .......... .......... .......... .......... 51% 2.36M 3s
  1700K .......... .......... .......... .......... .......... 52%  611M 3s
  1750K .......... .......... .......... .......... .......... 54%  231M 3s
  1800K .......... .......... .......... .......... .......... 55% 2.62M 3s
  1850K .......... .......... .......... .......... .......... 57%  151M 3s
  1900K .......... .......... .......... .......... .......... 58% 2.95M 3s
  1950K .......... .......... .......... .......... .......... 60% 61.9M 2s
  2000K .......... .......... .......... .......... .......... 61%  110M 2s
  2050K .......... .......... .......... .......... .......... 63% 3.23M 2s
  2100K .......... .......... .......... .......... .......... 65% 71.2M 2s
  2150K .......... .......... .......... .......... .......... 66% 72.1M 2s
  2200K .......... .......... .......... .......... .......... 68% 3.28M 2s
  2250K .......... .......... .......... .......... .......... 69% 66.7M 2s
  2300K .......... .......... .......... .......... .......... 71% 56.2M 2s
  2350K .......... .......... .......... .......... .......... 72% 3.40M 2s
  2400K .......... .......... .......... .......... .......... 74% 49.4M 1s
  2450K .......... .......... .......... .......... .......... 75% 51.8M 1s
  2500K .......... .......... .......... .......... .......... 77% 3.42M 1s
  2550K .......... .......... .......... .......... .......... 78% 52.0M 1s
  2600K .......... .......... .......... .......... .......... 80% 55.0M 1s
  2650K .......... .......... .......... .......... .......... 81% 3.40M 1s
  2700K .......... .......... .......... .......... .......... 83% 88.0M 1s
  2750K .......... .......... .......... .......... .......... 84% 49.0M 1s
  2800K .......... .......... .......... .......... .......... 86% 3.41M 1s
  2850K .......... .......... .......... .......... .......... 87% 74.1M 1s
  2900K .......... .......... .......... .......... .......... 89% 54.9M 1s
  2950K .......... .......... .......... .......... .......... 90% 4.67M 0s
  3000K .......... .......... .......... .......... .......... 92% 10.7M 0s
  3050K .......... .......... .......... .......... .......... 93%  103M 0s
  3100K .......... .......... .......... .......... .......... 95% 41.4M 0s
  3150K .......... .......... .......... .......... .......... 96% 3.50M 0s
  3200K .......... .......... .......... .......... .......... 98% 72.1M 0s
  3250K .......... .......... .......... .......... .......... 99% 93.5M 0s
  3300K ......                                                100% 42.8M=4.8s

2020-03-02 03:24:13 (5.61 Mb/s) - ‘/dev/null’ saved [3385841/3385841]

