--2020-03-02 03:23:45--  http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D419
Resolving biblioteca.inu.edu.sv (biblioteca.inu.edu.sv)... 78.47.62.221
Connecting to biblioteca.inu.edu.sv (biblioteca.inu.edu.sv)|78.47.62.221|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D419/ [following]
--2020-03-02 03:23:46--  http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D419/
Reusing existing connection to biblioteca.inu.edu.sv:80.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 3.22M
    50K .......... .......... .......... .......... .......... 5.14M
   100K .......... ....                                        26.1M=0.2s

2020-03-02 03:23:46 (4.44 Mb/s) - ‘/dev/null’ saved [117462]

--2020-03-02 03:23:46--  http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D387
Resolving biblioteca.inu.edu.sv (biblioteca.inu.edu.sv)... 78.47.62.221
Connecting to biblioteca.inu.edu.sv (biblioteca.inu.edu.sv)|78.47.62.221|:80... connected.
HTTP request sent, awaiting response... 301 Moved Permanently
Location: http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D387/ [following]
--2020-03-02 03:23:46--  http://biblioteca.inu.edu.sv/%3Fwpfb_dl%3D387/
Reusing existing connection to biblioteca.inu.edu.sv:80.
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 3.37M
    50K .......... .......... .......... .......... .......... 3.16M
   100K .......... ....                                        25.8M=0.3s

2020-03-02 03:23:47 (3.68 Mb/s) - ‘/dev/null’ saved [117462]

