--2020-03-02 03:24:16--  http://www.tsc.gob.sv/pdf/constitucionsv.pdf
Resolving www.tsc.gob.sv (www.tsc.gob.sv)... 104.27.170.247, 104.27.171.247
Connecting to www.tsc.gob.sv (www.tsc.gob.sv)|104.27.170.247|:80... connected.
HTTP request sent, awaiting response... 200 OK
Length: 249063 (243K) [application/pdf]
Saving to: ‘/dev/null’

     0K .......... .......... .......... .......... .......... 20% 34.8M 0s
    50K .......... .......... .......... .......... .......... 41% 5.00M 0s
   100K .......... .......... .......... .......... .......... 61% 80.8M 0s
   150K .......... .......... .......... .......... .......... 82% 5.33M 0s
   200K .......... .......... .......... .......... ...       100% 96.0M=0.2s

2020-03-02 03:24:17 (11.1 Mb/s) - ‘/dev/null’ saved [249063/249063]

