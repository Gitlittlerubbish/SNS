--2020-02-25 22:12:59--  http://www.upan.edu.sv/pdf/catalogo2017.pdf%0D
Resolving www.upan.edu.sv (www.upan.edu.sv)... 143.95.150.52
Connecting to www.upan.edu.sv (www.upan.edu.sv)|143.95.150.52|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:01 ERROR 404: Not Found.

--2020-02-25 22:13:34--  http://www.upan.edu.sv/pdf/catalogo2017.pdf%0D
Resolving www.upan.edu.sv (www.upan.edu.sv)... 143.95.150.52
Connecting to www.upan.edu.sv (www.upan.edu.sv)|143.95.150.52|:80... connected.
HTTP request sent, awaiting response... 404 Not Found
2020-02-25 22:13:35 ERROR 404: Not Found.

